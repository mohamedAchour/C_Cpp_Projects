// core.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module core (
		input  wire        clk_clk,                         //    clk.clk
		output wire        hps_io_hps_io_emac1_inst_TX_CLK, // hps_io.hps_io_emac1_inst_TX_CLK
		output wire        hps_io_hps_io_emac1_inst_TXD0,   //       .hps_io_emac1_inst_TXD0
		output wire        hps_io_hps_io_emac1_inst_TXD1,   //       .hps_io_emac1_inst_TXD1
		output wire        hps_io_hps_io_emac1_inst_TXD2,   //       .hps_io_emac1_inst_TXD2
		output wire        hps_io_hps_io_emac1_inst_TXD3,   //       .hps_io_emac1_inst_TXD3
		input  wire        hps_io_hps_io_emac1_inst_RXD0,   //       .hps_io_emac1_inst_RXD0
		inout  wire        hps_io_hps_io_emac1_inst_MDIO,   //       .hps_io_emac1_inst_MDIO
		output wire        hps_io_hps_io_emac1_inst_MDC,    //       .hps_io_emac1_inst_MDC
		input  wire        hps_io_hps_io_emac1_inst_RX_CTL, //       .hps_io_emac1_inst_RX_CTL
		output wire        hps_io_hps_io_emac1_inst_TX_CTL, //       .hps_io_emac1_inst_TX_CTL
		input  wire        hps_io_hps_io_emac1_inst_RX_CLK, //       .hps_io_emac1_inst_RX_CLK
		input  wire        hps_io_hps_io_emac1_inst_RXD1,   //       .hps_io_emac1_inst_RXD1
		input  wire        hps_io_hps_io_emac1_inst_RXD2,   //       .hps_io_emac1_inst_RXD2
		input  wire        hps_io_hps_io_emac1_inst_RXD3,   //       .hps_io_emac1_inst_RXD3
		inout  wire        hps_io_hps_io_sdio_inst_CMD,     //       .hps_io_sdio_inst_CMD
		inout  wire        hps_io_hps_io_sdio_inst_D0,      //       .hps_io_sdio_inst_D0
		inout  wire        hps_io_hps_io_sdio_inst_D1,      //       .hps_io_sdio_inst_D1
		output wire        hps_io_hps_io_sdio_inst_CLK,     //       .hps_io_sdio_inst_CLK
		inout  wire        hps_io_hps_io_sdio_inst_D2,      //       .hps_io_sdio_inst_D2
		inout  wire        hps_io_hps_io_sdio_inst_D3,      //       .hps_io_sdio_inst_D3
		input  wire        hps_io_hps_io_uart0_inst_RX,     //       .hps_io_uart0_inst_RX
		output wire        hps_io_hps_io_uart0_inst_TX,     //       .hps_io_uart0_inst_TX
		inout  wire        hps_io_hps_io_i2c0_inst_SDA,     //       .hps_io_i2c0_inst_SDA
		inout  wire        hps_io_hps_io_i2c0_inst_SCL,     //       .hps_io_i2c0_inst_SCL
		inout  wire        hps_io_hps_io_i2c1_inst_SDA,     //       .hps_io_i2c1_inst_SDA
		inout  wire        hps_io_hps_io_i2c1_inst_SCL,     //       .hps_io_i2c1_inst_SCL
		output wire [14:0] memory_mem_a,                    // memory.mem_a
		output wire [2:0]  memory_mem_ba,                   //       .mem_ba
		output wire        memory_mem_ck,                   //       .mem_ck
		output wire        memory_mem_ck_n,                 //       .mem_ck_n
		output wire        memory_mem_cke,                  //       .mem_cke
		output wire        memory_mem_cs_n,                 //       .mem_cs_n
		output wire        memory_mem_ras_n,                //       .mem_ras_n
		output wire        memory_mem_cas_n,                //       .mem_cas_n
		output wire        memory_mem_we_n,                 //       .mem_we_n
		output wire        memory_mem_reset_n,              //       .mem_reset_n
		inout  wire [31:0] memory_mem_dq,                   //       .mem_dq
		inout  wire [3:0]  memory_mem_dqs,                  //       .mem_dqs
		inout  wire [3:0]  memory_mem_dqs_n,                //       .mem_dqs_n
		output wire        memory_mem_odt,                  //       .mem_odt
		output wire [3:0]  memory_mem_dm,                   //       .mem_dm
		input  wire        memory_oct_rzqin,                //       .oct_rzqin
		output wire        pwm_a_pwm,                       //    pwm.a_pwm
		output wire        pwm_b_pwm,                       //       .b_pwm
		input  wire        pwm_secure,                      //       .secure
		input  wire        reset_reset_n                    //  reset.reset_n
	);

	wire         pll_0_outclk0_clk;                                                  // pll_0:outclk_0 -> [a_4_quadrant_chopper_0:csi_clock, mm_interconnect_0:pll_0_outclk0_clk, rst_controller:clk]
	wire   [1:0] hps_system_h2f_lw_axi_master_awburst;                               // hps_system:h2f_lw_AWBURST -> mm_interconnect_0:hps_system_h2f_lw_axi_master_awburst
	wire   [3:0] hps_system_h2f_lw_axi_master_arlen;                                 // hps_system:h2f_lw_ARLEN -> mm_interconnect_0:hps_system_h2f_lw_axi_master_arlen
	wire   [3:0] hps_system_h2f_lw_axi_master_wstrb;                                 // hps_system:h2f_lw_WSTRB -> mm_interconnect_0:hps_system_h2f_lw_axi_master_wstrb
	wire         hps_system_h2f_lw_axi_master_wready;                                // mm_interconnect_0:hps_system_h2f_lw_axi_master_wready -> hps_system:h2f_lw_WREADY
	wire  [11:0] hps_system_h2f_lw_axi_master_rid;                                   // mm_interconnect_0:hps_system_h2f_lw_axi_master_rid -> hps_system:h2f_lw_RID
	wire         hps_system_h2f_lw_axi_master_rready;                                // hps_system:h2f_lw_RREADY -> mm_interconnect_0:hps_system_h2f_lw_axi_master_rready
	wire   [3:0] hps_system_h2f_lw_axi_master_awlen;                                 // hps_system:h2f_lw_AWLEN -> mm_interconnect_0:hps_system_h2f_lw_axi_master_awlen
	wire  [11:0] hps_system_h2f_lw_axi_master_wid;                                   // hps_system:h2f_lw_WID -> mm_interconnect_0:hps_system_h2f_lw_axi_master_wid
	wire   [3:0] hps_system_h2f_lw_axi_master_arcache;                               // hps_system:h2f_lw_ARCACHE -> mm_interconnect_0:hps_system_h2f_lw_axi_master_arcache
	wire         hps_system_h2f_lw_axi_master_wvalid;                                // hps_system:h2f_lw_WVALID -> mm_interconnect_0:hps_system_h2f_lw_axi_master_wvalid
	wire  [20:0] hps_system_h2f_lw_axi_master_araddr;                                // hps_system:h2f_lw_ARADDR -> mm_interconnect_0:hps_system_h2f_lw_axi_master_araddr
	wire   [2:0] hps_system_h2f_lw_axi_master_arprot;                                // hps_system:h2f_lw_ARPROT -> mm_interconnect_0:hps_system_h2f_lw_axi_master_arprot
	wire   [2:0] hps_system_h2f_lw_axi_master_awprot;                                // hps_system:h2f_lw_AWPROT -> mm_interconnect_0:hps_system_h2f_lw_axi_master_awprot
	wire  [31:0] hps_system_h2f_lw_axi_master_wdata;                                 // hps_system:h2f_lw_WDATA -> mm_interconnect_0:hps_system_h2f_lw_axi_master_wdata
	wire         hps_system_h2f_lw_axi_master_arvalid;                               // hps_system:h2f_lw_ARVALID -> mm_interconnect_0:hps_system_h2f_lw_axi_master_arvalid
	wire   [3:0] hps_system_h2f_lw_axi_master_awcache;                               // hps_system:h2f_lw_AWCACHE -> mm_interconnect_0:hps_system_h2f_lw_axi_master_awcache
	wire  [11:0] hps_system_h2f_lw_axi_master_arid;                                  // hps_system:h2f_lw_ARID -> mm_interconnect_0:hps_system_h2f_lw_axi_master_arid
	wire   [1:0] hps_system_h2f_lw_axi_master_arlock;                                // hps_system:h2f_lw_ARLOCK -> mm_interconnect_0:hps_system_h2f_lw_axi_master_arlock
	wire   [1:0] hps_system_h2f_lw_axi_master_awlock;                                // hps_system:h2f_lw_AWLOCK -> mm_interconnect_0:hps_system_h2f_lw_axi_master_awlock
	wire  [20:0] hps_system_h2f_lw_axi_master_awaddr;                                // hps_system:h2f_lw_AWADDR -> mm_interconnect_0:hps_system_h2f_lw_axi_master_awaddr
	wire   [1:0] hps_system_h2f_lw_axi_master_bresp;                                 // mm_interconnect_0:hps_system_h2f_lw_axi_master_bresp -> hps_system:h2f_lw_BRESP
	wire         hps_system_h2f_lw_axi_master_arready;                               // mm_interconnect_0:hps_system_h2f_lw_axi_master_arready -> hps_system:h2f_lw_ARREADY
	wire  [31:0] hps_system_h2f_lw_axi_master_rdata;                                 // mm_interconnect_0:hps_system_h2f_lw_axi_master_rdata -> hps_system:h2f_lw_RDATA
	wire         hps_system_h2f_lw_axi_master_awready;                               // mm_interconnect_0:hps_system_h2f_lw_axi_master_awready -> hps_system:h2f_lw_AWREADY
	wire   [1:0] hps_system_h2f_lw_axi_master_arburst;                               // hps_system:h2f_lw_ARBURST -> mm_interconnect_0:hps_system_h2f_lw_axi_master_arburst
	wire   [2:0] hps_system_h2f_lw_axi_master_arsize;                                // hps_system:h2f_lw_ARSIZE -> mm_interconnect_0:hps_system_h2f_lw_axi_master_arsize
	wire         hps_system_h2f_lw_axi_master_bready;                                // hps_system:h2f_lw_BREADY -> mm_interconnect_0:hps_system_h2f_lw_axi_master_bready
	wire         hps_system_h2f_lw_axi_master_rlast;                                 // mm_interconnect_0:hps_system_h2f_lw_axi_master_rlast -> hps_system:h2f_lw_RLAST
	wire         hps_system_h2f_lw_axi_master_wlast;                                 // hps_system:h2f_lw_WLAST -> mm_interconnect_0:hps_system_h2f_lw_axi_master_wlast
	wire   [1:0] hps_system_h2f_lw_axi_master_rresp;                                 // mm_interconnect_0:hps_system_h2f_lw_axi_master_rresp -> hps_system:h2f_lw_RRESP
	wire  [11:0] hps_system_h2f_lw_axi_master_awid;                                  // hps_system:h2f_lw_AWID -> mm_interconnect_0:hps_system_h2f_lw_axi_master_awid
	wire  [11:0] hps_system_h2f_lw_axi_master_bid;                                   // mm_interconnect_0:hps_system_h2f_lw_axi_master_bid -> hps_system:h2f_lw_BID
	wire         hps_system_h2f_lw_axi_master_bvalid;                                // mm_interconnect_0:hps_system_h2f_lw_axi_master_bvalid -> hps_system:h2f_lw_BVALID
	wire   [2:0] hps_system_h2f_lw_axi_master_awsize;                                // hps_system:h2f_lw_AWSIZE -> mm_interconnect_0:hps_system_h2f_lw_axi_master_awsize
	wire         hps_system_h2f_lw_axi_master_awvalid;                               // hps_system:h2f_lw_AWVALID -> mm_interconnect_0:hps_system_h2f_lw_axi_master_awvalid
	wire         hps_system_h2f_lw_axi_master_rvalid;                                // mm_interconnect_0:hps_system_h2f_lw_axi_master_rvalid -> hps_system:h2f_lw_RVALID
	wire  [31:0] master_jtag_master_readdata;                                        // mm_interconnect_0:master_jtag_master_readdata -> master_jtag:master_readdata
	wire         master_jtag_master_waitrequest;                                     // mm_interconnect_0:master_jtag_master_waitrequest -> master_jtag:master_waitrequest
	wire  [31:0] master_jtag_master_address;                                         // master_jtag:master_address -> mm_interconnect_0:master_jtag_master_address
	wire         master_jtag_master_read;                                            // master_jtag:master_read -> mm_interconnect_0:master_jtag_master_read
	wire   [3:0] master_jtag_master_byteenable;                                      // master_jtag:master_byteenable -> mm_interconnect_0:master_jtag_master_byteenable
	wire         master_jtag_master_readdatavalid;                                   // mm_interconnect_0:master_jtag_master_readdatavalid -> master_jtag:master_readdatavalid
	wire         master_jtag_master_write;                                           // master_jtag:master_write -> mm_interconnect_0:master_jtag_master_write
	wire  [31:0] master_jtag_master_writedata;                                       // master_jtag:master_writedata -> mm_interconnect_0:master_jtag_master_writedata
	wire  [15:0] mm_interconnect_0_a_4_quadrant_chopper_0_avalon_slave_0_readdata;   // a_4_quadrant_chopper_0:avs_readdata -> mm_interconnect_0:a_4_quadrant_chopper_0_avalon_slave_0_readdata
	wire   [1:0] mm_interconnect_0_a_4_quadrant_chopper_0_avalon_slave_0_address;    // mm_interconnect_0:a_4_quadrant_chopper_0_avalon_slave_0_address -> a_4_quadrant_chopper_0:avs_address
	wire         mm_interconnect_0_a_4_quadrant_chopper_0_avalon_slave_0_read;       // mm_interconnect_0:a_4_quadrant_chopper_0_avalon_slave_0_read -> a_4_quadrant_chopper_0:avs_read
	wire   [1:0] mm_interconnect_0_a_4_quadrant_chopper_0_avalon_slave_0_byteenable; // mm_interconnect_0:a_4_quadrant_chopper_0_avalon_slave_0_byteenable -> a_4_quadrant_chopper_0:avs_byteenable
	wire         mm_interconnect_0_a_4_quadrant_chopper_0_avalon_slave_0_write;      // mm_interconnect_0:a_4_quadrant_chopper_0_avalon_slave_0_write -> a_4_quadrant_chopper_0:avs_write
	wire  [15:0] mm_interconnect_0_a_4_quadrant_chopper_0_avalon_slave_0_writedata;  // mm_interconnect_0:a_4_quadrant_chopper_0_avalon_slave_0_writedata -> a_4_quadrant_chopper_0:avs_writedata
	wire  [31:0] mm_interconnect_0_sysid_control_slave_readdata;                     // sysid:readdata -> mm_interconnect_0:sysid_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_control_slave_address;                      // mm_interconnect_0:sysid_control_slave_address -> sysid:address
	wire         irq_mapper_receiver0_irq;                                           // a_4_quadrant_chopper_0:ins_end_cycle -> irq_mapper:receiver0_irq
	wire  [31:0] hps_system_f2h_irq0_irq;                                            // irq_mapper:sender_irq -> hps_system:f2h_irq_p0
	wire  [31:0] hps_system_f2h_irq1_irq;                                            // irq_mapper_001:sender_irq -> hps_system:f2h_irq_p1
	wire         rst_controller_reset_out_reset;                                     // rst_controller:reset_out -> [a_4_quadrant_chopper_0:rsi_reset, mm_interconnect_0:a_4_quadrant_chopper_0_clock_reset_reset_bridge_in_reset_reset]
	wire         rst_controller_001_reset_out_reset;                                 // rst_controller_001:reset_out -> [mm_interconnect_0:master_jtag_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_0:sysid_reset_reset_bridge_in_reset_reset, sysid:reset_n]
	wire         rst_controller_002_reset_out_reset;                                 // rst_controller_002:reset_out -> mm_interconnect_0:hps_system_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset
	wire         hps_system_h2f_reset_reset;                                         // hps_system:h2f_rst_n -> rst_controller_002:reset_in0

	hacheur_top a_4_quadrant_chopper_0 (
		.rsi_reset      (rst_controller_reset_out_reset),                                     //        clock_reset.reset
		.avs_address    (mm_interconnect_0_a_4_quadrant_chopper_0_avalon_slave_0_address),    //     avalon_slave_0.address
		.avs_byteenable (mm_interconnect_0_a_4_quadrant_chopper_0_avalon_slave_0_byteenable), //                   .byteenable
		.avs_read       (mm_interconnect_0_a_4_quadrant_chopper_0_avalon_slave_0_read),       //                   .read
		.avs_readdata   (mm_interconnect_0_a_4_quadrant_chopper_0_avalon_slave_0_readdata),   //                   .readdata
		.avs_write      (mm_interconnect_0_a_4_quadrant_chopper_0_avalon_slave_0_write),      //                   .write
		.avs_writedata  (mm_interconnect_0_a_4_quadrant_chopper_0_avalon_slave_0_writedata),  //                   .writedata
		.ins_end_cycle  (irq_mapper_receiver0_irq),                                           // interrupt_sender_0.irq_n
		.csi_clock      (pll_0_outclk0_clk),                                                  //         clock_sink.clk
		.A              (pwm_a_pwm),                                                          //        conduit_end.a_pwm
		.B              (pwm_b_pwm),                                                          //                   .b_pwm
		.secure         (pwm_secure)                                                          //                   .secure
	);

	core_hps_system #(
		.F2S_Width (2),
		.S2F_Width (2)
	) hps_system (
		.h2f_mpu_eventi           (),                                     //    h2f_mpu_events.eventi
		.h2f_mpu_evento           (),                                     //                  .evento
		.h2f_mpu_standbywfe       (),                                     //                  .standbywfe
		.h2f_mpu_standbywfi       (),                                     //                  .standbywfi
		.mem_a                    (memory_mem_a),                         //            memory.mem_a
		.mem_ba                   (memory_mem_ba),                        //                  .mem_ba
		.mem_ck                   (memory_mem_ck),                        //                  .mem_ck
		.mem_ck_n                 (memory_mem_ck_n),                      //                  .mem_ck_n
		.mem_cke                  (memory_mem_cke),                       //                  .mem_cke
		.mem_cs_n                 (memory_mem_cs_n),                      //                  .mem_cs_n
		.mem_ras_n                (memory_mem_ras_n),                     //                  .mem_ras_n
		.mem_cas_n                (memory_mem_cas_n),                     //                  .mem_cas_n
		.mem_we_n                 (memory_mem_we_n),                      //                  .mem_we_n
		.mem_reset_n              (memory_mem_reset_n),                   //                  .mem_reset_n
		.mem_dq                   (memory_mem_dq),                        //                  .mem_dq
		.mem_dqs                  (memory_mem_dqs),                       //                  .mem_dqs
		.mem_dqs_n                (memory_mem_dqs_n),                     //                  .mem_dqs_n
		.mem_odt                  (memory_mem_odt),                       //                  .mem_odt
		.mem_dm                   (memory_mem_dm),                        //                  .mem_dm
		.oct_rzqin                (memory_oct_rzqin),                     //                  .oct_rzqin
		.hps_io_emac1_inst_TX_CLK (hps_io_hps_io_emac1_inst_TX_CLK),      //            hps_io.hps_io_emac1_inst_TX_CLK
		.hps_io_emac1_inst_TXD0   (hps_io_hps_io_emac1_inst_TXD0),        //                  .hps_io_emac1_inst_TXD0
		.hps_io_emac1_inst_TXD1   (hps_io_hps_io_emac1_inst_TXD1),        //                  .hps_io_emac1_inst_TXD1
		.hps_io_emac1_inst_TXD2   (hps_io_hps_io_emac1_inst_TXD2),        //                  .hps_io_emac1_inst_TXD2
		.hps_io_emac1_inst_TXD3   (hps_io_hps_io_emac1_inst_TXD3),        //                  .hps_io_emac1_inst_TXD3
		.hps_io_emac1_inst_RXD0   (hps_io_hps_io_emac1_inst_RXD0),        //                  .hps_io_emac1_inst_RXD0
		.hps_io_emac1_inst_MDIO   (hps_io_hps_io_emac1_inst_MDIO),        //                  .hps_io_emac1_inst_MDIO
		.hps_io_emac1_inst_MDC    (hps_io_hps_io_emac1_inst_MDC),         //                  .hps_io_emac1_inst_MDC
		.hps_io_emac1_inst_RX_CTL (hps_io_hps_io_emac1_inst_RX_CTL),      //                  .hps_io_emac1_inst_RX_CTL
		.hps_io_emac1_inst_TX_CTL (hps_io_hps_io_emac1_inst_TX_CTL),      //                  .hps_io_emac1_inst_TX_CTL
		.hps_io_emac1_inst_RX_CLK (hps_io_hps_io_emac1_inst_RX_CLK),      //                  .hps_io_emac1_inst_RX_CLK
		.hps_io_emac1_inst_RXD1   (hps_io_hps_io_emac1_inst_RXD1),        //                  .hps_io_emac1_inst_RXD1
		.hps_io_emac1_inst_RXD2   (hps_io_hps_io_emac1_inst_RXD2),        //                  .hps_io_emac1_inst_RXD2
		.hps_io_emac1_inst_RXD3   (hps_io_hps_io_emac1_inst_RXD3),        //                  .hps_io_emac1_inst_RXD3
		.hps_io_sdio_inst_CMD     (hps_io_hps_io_sdio_inst_CMD),          //                  .hps_io_sdio_inst_CMD
		.hps_io_sdio_inst_D0      (hps_io_hps_io_sdio_inst_D0),           //                  .hps_io_sdio_inst_D0
		.hps_io_sdio_inst_D1      (hps_io_hps_io_sdio_inst_D1),           //                  .hps_io_sdio_inst_D1
		.hps_io_sdio_inst_CLK     (hps_io_hps_io_sdio_inst_CLK),          //                  .hps_io_sdio_inst_CLK
		.hps_io_sdio_inst_D2      (hps_io_hps_io_sdio_inst_D2),           //                  .hps_io_sdio_inst_D2
		.hps_io_sdio_inst_D3      (hps_io_hps_io_sdio_inst_D3),           //                  .hps_io_sdio_inst_D3
		.hps_io_uart0_inst_RX     (hps_io_hps_io_uart0_inst_RX),          //                  .hps_io_uart0_inst_RX
		.hps_io_uart0_inst_TX     (hps_io_hps_io_uart0_inst_TX),          //                  .hps_io_uart0_inst_TX
		.hps_io_i2c0_inst_SDA     (hps_io_hps_io_i2c0_inst_SDA),          //                  .hps_io_i2c0_inst_SDA
		.hps_io_i2c0_inst_SCL     (hps_io_hps_io_i2c0_inst_SCL),          //                  .hps_io_i2c0_inst_SCL
		.hps_io_i2c1_inst_SDA     (hps_io_hps_io_i2c1_inst_SDA),          //                  .hps_io_i2c1_inst_SDA
		.hps_io_i2c1_inst_SCL     (hps_io_hps_io_i2c1_inst_SCL),          //                  .hps_io_i2c1_inst_SCL
		.h2f_rst_n                (hps_system_h2f_reset_reset),           //         h2f_reset.reset_n
		.f2h_sdram0_clk           (clk_clk),                              //  f2h_sdram0_clock.clk
		.f2h_sdram0_ARADDR        (),                                     //   f2h_sdram0_data.araddr
		.f2h_sdram0_ARLEN         (),                                     //                  .arlen
		.f2h_sdram0_ARID          (),                                     //                  .arid
		.f2h_sdram0_ARSIZE        (),                                     //                  .arsize
		.f2h_sdram0_ARBURST       (),                                     //                  .arburst
		.f2h_sdram0_ARLOCK        (),                                     //                  .arlock
		.f2h_sdram0_ARPROT        (),                                     //                  .arprot
		.f2h_sdram0_ARVALID       (),                                     //                  .arvalid
		.f2h_sdram0_ARCACHE       (),                                     //                  .arcache
		.f2h_sdram0_AWADDR        (),                                     //                  .awaddr
		.f2h_sdram0_AWLEN         (),                                     //                  .awlen
		.f2h_sdram0_AWID          (),                                     //                  .awid
		.f2h_sdram0_AWSIZE        (),                                     //                  .awsize
		.f2h_sdram0_AWBURST       (),                                     //                  .awburst
		.f2h_sdram0_AWLOCK        (),                                     //                  .awlock
		.f2h_sdram0_AWPROT        (),                                     //                  .awprot
		.f2h_sdram0_AWVALID       (),                                     //                  .awvalid
		.f2h_sdram0_AWCACHE       (),                                     //                  .awcache
		.f2h_sdram0_BRESP         (),                                     //                  .bresp
		.f2h_sdram0_BID           (),                                     //                  .bid
		.f2h_sdram0_BVALID        (),                                     //                  .bvalid
		.f2h_sdram0_BREADY        (),                                     //                  .bready
		.f2h_sdram0_ARREADY       (),                                     //                  .arready
		.f2h_sdram0_AWREADY       (),                                     //                  .awready
		.f2h_sdram0_RREADY        (),                                     //                  .rready
		.f2h_sdram0_RDATA         (),                                     //                  .rdata
		.f2h_sdram0_RRESP         (),                                     //                  .rresp
		.f2h_sdram0_RLAST         (),                                     //                  .rlast
		.f2h_sdram0_RID           (),                                     //                  .rid
		.f2h_sdram0_RVALID        (),                                     //                  .rvalid
		.f2h_sdram0_WLAST         (),                                     //                  .wlast
		.f2h_sdram0_WVALID        (),                                     //                  .wvalid
		.f2h_sdram0_WDATA         (),                                     //                  .wdata
		.f2h_sdram0_WSTRB         (),                                     //                  .wstrb
		.f2h_sdram0_WREADY        (),                                     //                  .wready
		.f2h_sdram0_WID           (),                                     //                  .wid
		.h2f_axi_clk              (clk_clk),                              //     h2f_axi_clock.clk
		.h2f_AWID                 (),                                     //    h2f_axi_master.awid
		.h2f_AWADDR               (),                                     //                  .awaddr
		.h2f_AWLEN                (),                                     //                  .awlen
		.h2f_AWSIZE               (),                                     //                  .awsize
		.h2f_AWBURST              (),                                     //                  .awburst
		.h2f_AWLOCK               (),                                     //                  .awlock
		.h2f_AWCACHE              (),                                     //                  .awcache
		.h2f_AWPROT               (),                                     //                  .awprot
		.h2f_AWVALID              (),                                     //                  .awvalid
		.h2f_AWREADY              (),                                     //                  .awready
		.h2f_WID                  (),                                     //                  .wid
		.h2f_WDATA                (),                                     //                  .wdata
		.h2f_WSTRB                (),                                     //                  .wstrb
		.h2f_WLAST                (),                                     //                  .wlast
		.h2f_WVALID               (),                                     //                  .wvalid
		.h2f_WREADY               (),                                     //                  .wready
		.h2f_BID                  (),                                     //                  .bid
		.h2f_BRESP                (),                                     //                  .bresp
		.h2f_BVALID               (),                                     //                  .bvalid
		.h2f_BREADY               (),                                     //                  .bready
		.h2f_ARID                 (),                                     //                  .arid
		.h2f_ARADDR               (),                                     //                  .araddr
		.h2f_ARLEN                (),                                     //                  .arlen
		.h2f_ARSIZE               (),                                     //                  .arsize
		.h2f_ARBURST              (),                                     //                  .arburst
		.h2f_ARLOCK               (),                                     //                  .arlock
		.h2f_ARCACHE              (),                                     //                  .arcache
		.h2f_ARPROT               (),                                     //                  .arprot
		.h2f_ARVALID              (),                                     //                  .arvalid
		.h2f_ARREADY              (),                                     //                  .arready
		.h2f_RID                  (),                                     //                  .rid
		.h2f_RDATA                (),                                     //                  .rdata
		.h2f_RRESP                (),                                     //                  .rresp
		.h2f_RLAST                (),                                     //                  .rlast
		.h2f_RVALID               (),                                     //                  .rvalid
		.h2f_RREADY               (),                                     //                  .rready
		.f2h_axi_clk              (clk_clk),                              //     f2h_axi_clock.clk
		.f2h_AWID                 (),                                     //     f2h_axi_slave.awid
		.f2h_AWADDR               (),                                     //                  .awaddr
		.f2h_AWLEN                (),                                     //                  .awlen
		.f2h_AWSIZE               (),                                     //                  .awsize
		.f2h_AWBURST              (),                                     //                  .awburst
		.f2h_AWLOCK               (),                                     //                  .awlock
		.f2h_AWCACHE              (),                                     //                  .awcache
		.f2h_AWPROT               (),                                     //                  .awprot
		.f2h_AWVALID              (),                                     //                  .awvalid
		.f2h_AWREADY              (),                                     //                  .awready
		.f2h_AWUSER               (),                                     //                  .awuser
		.f2h_WID                  (),                                     //                  .wid
		.f2h_WDATA                (),                                     //                  .wdata
		.f2h_WSTRB                (),                                     //                  .wstrb
		.f2h_WLAST                (),                                     //                  .wlast
		.f2h_WVALID               (),                                     //                  .wvalid
		.f2h_WREADY               (),                                     //                  .wready
		.f2h_BID                  (),                                     //                  .bid
		.f2h_BRESP                (),                                     //                  .bresp
		.f2h_BVALID               (),                                     //                  .bvalid
		.f2h_BREADY               (),                                     //                  .bready
		.f2h_ARID                 (),                                     //                  .arid
		.f2h_ARADDR               (),                                     //                  .araddr
		.f2h_ARLEN                (),                                     //                  .arlen
		.f2h_ARSIZE               (),                                     //                  .arsize
		.f2h_ARBURST              (),                                     //                  .arburst
		.f2h_ARLOCK               (),                                     //                  .arlock
		.f2h_ARCACHE              (),                                     //                  .arcache
		.f2h_ARPROT               (),                                     //                  .arprot
		.f2h_ARVALID              (),                                     //                  .arvalid
		.f2h_ARREADY              (),                                     //                  .arready
		.f2h_ARUSER               (),                                     //                  .aruser
		.f2h_RID                  (),                                     //                  .rid
		.f2h_RDATA                (),                                     //                  .rdata
		.f2h_RRESP                (),                                     //                  .rresp
		.f2h_RLAST                (),                                     //                  .rlast
		.f2h_RVALID               (),                                     //                  .rvalid
		.f2h_RREADY               (),                                     //                  .rready
		.h2f_lw_axi_clk           (clk_clk),                              //  h2f_lw_axi_clock.clk
		.h2f_lw_AWID              (hps_system_h2f_lw_axi_master_awid),    // h2f_lw_axi_master.awid
		.h2f_lw_AWADDR            (hps_system_h2f_lw_axi_master_awaddr),  //                  .awaddr
		.h2f_lw_AWLEN             (hps_system_h2f_lw_axi_master_awlen),   //                  .awlen
		.h2f_lw_AWSIZE            (hps_system_h2f_lw_axi_master_awsize),  //                  .awsize
		.h2f_lw_AWBURST           (hps_system_h2f_lw_axi_master_awburst), //                  .awburst
		.h2f_lw_AWLOCK            (hps_system_h2f_lw_axi_master_awlock),  //                  .awlock
		.h2f_lw_AWCACHE           (hps_system_h2f_lw_axi_master_awcache), //                  .awcache
		.h2f_lw_AWPROT            (hps_system_h2f_lw_axi_master_awprot),  //                  .awprot
		.h2f_lw_AWVALID           (hps_system_h2f_lw_axi_master_awvalid), //                  .awvalid
		.h2f_lw_AWREADY           (hps_system_h2f_lw_axi_master_awready), //                  .awready
		.h2f_lw_WID               (hps_system_h2f_lw_axi_master_wid),     //                  .wid
		.h2f_lw_WDATA             (hps_system_h2f_lw_axi_master_wdata),   //                  .wdata
		.h2f_lw_WSTRB             (hps_system_h2f_lw_axi_master_wstrb),   //                  .wstrb
		.h2f_lw_WLAST             (hps_system_h2f_lw_axi_master_wlast),   //                  .wlast
		.h2f_lw_WVALID            (hps_system_h2f_lw_axi_master_wvalid),  //                  .wvalid
		.h2f_lw_WREADY            (hps_system_h2f_lw_axi_master_wready),  //                  .wready
		.h2f_lw_BID               (hps_system_h2f_lw_axi_master_bid),     //                  .bid
		.h2f_lw_BRESP             (hps_system_h2f_lw_axi_master_bresp),   //                  .bresp
		.h2f_lw_BVALID            (hps_system_h2f_lw_axi_master_bvalid),  //                  .bvalid
		.h2f_lw_BREADY            (hps_system_h2f_lw_axi_master_bready),  //                  .bready
		.h2f_lw_ARID              (hps_system_h2f_lw_axi_master_arid),    //                  .arid
		.h2f_lw_ARADDR            (hps_system_h2f_lw_axi_master_araddr),  //                  .araddr
		.h2f_lw_ARLEN             (hps_system_h2f_lw_axi_master_arlen),   //                  .arlen
		.h2f_lw_ARSIZE            (hps_system_h2f_lw_axi_master_arsize),  //                  .arsize
		.h2f_lw_ARBURST           (hps_system_h2f_lw_axi_master_arburst), //                  .arburst
		.h2f_lw_ARLOCK            (hps_system_h2f_lw_axi_master_arlock),  //                  .arlock
		.h2f_lw_ARCACHE           (hps_system_h2f_lw_axi_master_arcache), //                  .arcache
		.h2f_lw_ARPROT            (hps_system_h2f_lw_axi_master_arprot),  //                  .arprot
		.h2f_lw_ARVALID           (hps_system_h2f_lw_axi_master_arvalid), //                  .arvalid
		.h2f_lw_ARREADY           (hps_system_h2f_lw_axi_master_arready), //                  .arready
		.h2f_lw_RID               (hps_system_h2f_lw_axi_master_rid),     //                  .rid
		.h2f_lw_RDATA             (hps_system_h2f_lw_axi_master_rdata),   //                  .rdata
		.h2f_lw_RRESP             (hps_system_h2f_lw_axi_master_rresp),   //                  .rresp
		.h2f_lw_RLAST             (hps_system_h2f_lw_axi_master_rlast),   //                  .rlast
		.h2f_lw_RVALID            (hps_system_h2f_lw_axi_master_rvalid),  //                  .rvalid
		.h2f_lw_RREADY            (hps_system_h2f_lw_axi_master_rready),  //                  .rready
		.f2h_irq_p0               (hps_system_f2h_irq0_irq),              //          f2h_irq0.irq
		.f2h_irq_p1               (hps_system_f2h_irq1_irq)               //          f2h_irq1.irq
	);

	core_master_jtag #(
		.USE_PLI     (0),
		.PLI_PORT    (50000),
		.FIFO_DEPTHS (2)
	) master_jtag (
		.clk_clk              (clk_clk),                          //          clk.clk
		.clk_reset_reset      (~reset_reset_n),                   //    clk_reset.reset
		.master_address       (master_jtag_master_address),       //       master.address
		.master_readdata      (master_jtag_master_readdata),      //             .readdata
		.master_read          (master_jtag_master_read),          //             .read
		.master_write         (master_jtag_master_write),         //             .write
		.master_writedata     (master_jtag_master_writedata),     //             .writedata
		.master_waitrequest   (master_jtag_master_waitrequest),   //             .waitrequest
		.master_readdatavalid (master_jtag_master_readdatavalid), //             .readdatavalid
		.master_byteenable    (master_jtag_master_byteenable),    //             .byteenable
		.master_reset_reset   ()                                  // master_reset.reset
	);

	core_pll_0 pll_0 (
		.refclk   (clk_clk),           //  refclk.clk
		.rst      (~reset_reset_n),    //   reset.reset
		.outclk_0 (pll_0_outclk0_clk), // outclk0.clk
		.locked   ()                   // (terminated)
	);

	core_sysid sysid (
		.clock    (clk_clk),                                        //           clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),            //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_control_slave_address)   //              .address
	);

	core_mm_interconnect_0 mm_interconnect_0 (
		.hps_system_h2f_lw_axi_master_awid                                        (hps_system_h2f_lw_axi_master_awid),                                  //                                       hps_system_h2f_lw_axi_master.awid
		.hps_system_h2f_lw_axi_master_awaddr                                      (hps_system_h2f_lw_axi_master_awaddr),                                //                                                                   .awaddr
		.hps_system_h2f_lw_axi_master_awlen                                       (hps_system_h2f_lw_axi_master_awlen),                                 //                                                                   .awlen
		.hps_system_h2f_lw_axi_master_awsize                                      (hps_system_h2f_lw_axi_master_awsize),                                //                                                                   .awsize
		.hps_system_h2f_lw_axi_master_awburst                                     (hps_system_h2f_lw_axi_master_awburst),                               //                                                                   .awburst
		.hps_system_h2f_lw_axi_master_awlock                                      (hps_system_h2f_lw_axi_master_awlock),                                //                                                                   .awlock
		.hps_system_h2f_lw_axi_master_awcache                                     (hps_system_h2f_lw_axi_master_awcache),                               //                                                                   .awcache
		.hps_system_h2f_lw_axi_master_awprot                                      (hps_system_h2f_lw_axi_master_awprot),                                //                                                                   .awprot
		.hps_system_h2f_lw_axi_master_awvalid                                     (hps_system_h2f_lw_axi_master_awvalid),                               //                                                                   .awvalid
		.hps_system_h2f_lw_axi_master_awready                                     (hps_system_h2f_lw_axi_master_awready),                               //                                                                   .awready
		.hps_system_h2f_lw_axi_master_wid                                         (hps_system_h2f_lw_axi_master_wid),                                   //                                                                   .wid
		.hps_system_h2f_lw_axi_master_wdata                                       (hps_system_h2f_lw_axi_master_wdata),                                 //                                                                   .wdata
		.hps_system_h2f_lw_axi_master_wstrb                                       (hps_system_h2f_lw_axi_master_wstrb),                                 //                                                                   .wstrb
		.hps_system_h2f_lw_axi_master_wlast                                       (hps_system_h2f_lw_axi_master_wlast),                                 //                                                                   .wlast
		.hps_system_h2f_lw_axi_master_wvalid                                      (hps_system_h2f_lw_axi_master_wvalid),                                //                                                                   .wvalid
		.hps_system_h2f_lw_axi_master_wready                                      (hps_system_h2f_lw_axi_master_wready),                                //                                                                   .wready
		.hps_system_h2f_lw_axi_master_bid                                         (hps_system_h2f_lw_axi_master_bid),                                   //                                                                   .bid
		.hps_system_h2f_lw_axi_master_bresp                                       (hps_system_h2f_lw_axi_master_bresp),                                 //                                                                   .bresp
		.hps_system_h2f_lw_axi_master_bvalid                                      (hps_system_h2f_lw_axi_master_bvalid),                                //                                                                   .bvalid
		.hps_system_h2f_lw_axi_master_bready                                      (hps_system_h2f_lw_axi_master_bready),                                //                                                                   .bready
		.hps_system_h2f_lw_axi_master_arid                                        (hps_system_h2f_lw_axi_master_arid),                                  //                                                                   .arid
		.hps_system_h2f_lw_axi_master_araddr                                      (hps_system_h2f_lw_axi_master_araddr),                                //                                                                   .araddr
		.hps_system_h2f_lw_axi_master_arlen                                       (hps_system_h2f_lw_axi_master_arlen),                                 //                                                                   .arlen
		.hps_system_h2f_lw_axi_master_arsize                                      (hps_system_h2f_lw_axi_master_arsize),                                //                                                                   .arsize
		.hps_system_h2f_lw_axi_master_arburst                                     (hps_system_h2f_lw_axi_master_arburst),                               //                                                                   .arburst
		.hps_system_h2f_lw_axi_master_arlock                                      (hps_system_h2f_lw_axi_master_arlock),                                //                                                                   .arlock
		.hps_system_h2f_lw_axi_master_arcache                                     (hps_system_h2f_lw_axi_master_arcache),                               //                                                                   .arcache
		.hps_system_h2f_lw_axi_master_arprot                                      (hps_system_h2f_lw_axi_master_arprot),                                //                                                                   .arprot
		.hps_system_h2f_lw_axi_master_arvalid                                     (hps_system_h2f_lw_axi_master_arvalid),                               //                                                                   .arvalid
		.hps_system_h2f_lw_axi_master_arready                                     (hps_system_h2f_lw_axi_master_arready),                               //                                                                   .arready
		.hps_system_h2f_lw_axi_master_rid                                         (hps_system_h2f_lw_axi_master_rid),                                   //                                                                   .rid
		.hps_system_h2f_lw_axi_master_rdata                                       (hps_system_h2f_lw_axi_master_rdata),                                 //                                                                   .rdata
		.hps_system_h2f_lw_axi_master_rresp                                       (hps_system_h2f_lw_axi_master_rresp),                                 //                                                                   .rresp
		.hps_system_h2f_lw_axi_master_rlast                                       (hps_system_h2f_lw_axi_master_rlast),                                 //                                                                   .rlast
		.hps_system_h2f_lw_axi_master_rvalid                                      (hps_system_h2f_lw_axi_master_rvalid),                                //                                                                   .rvalid
		.hps_system_h2f_lw_axi_master_rready                                      (hps_system_h2f_lw_axi_master_rready),                                //                                                                   .rready
		.clk_0_clk_clk                                                            (clk_clk),                                                            //                                                          clk_0_clk.clk
		.pll_0_outclk0_clk                                                        (pll_0_outclk0_clk),                                                  //                                                      pll_0_outclk0.clk
		.a_4_quadrant_chopper_0_clock_reset_reset_bridge_in_reset_reset           (rst_controller_reset_out_reset),                                     //           a_4_quadrant_chopper_0_clock_reset_reset_bridge_in_reset.reset
		.hps_system_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset (rst_controller_002_reset_out_reset),                                 // hps_system_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
		.master_jtag_clk_reset_reset_bridge_in_reset_reset                        (rst_controller_001_reset_out_reset),                                 //                        master_jtag_clk_reset_reset_bridge_in_reset.reset
		.sysid_reset_reset_bridge_in_reset_reset                                  (rst_controller_001_reset_out_reset),                                 //                                  sysid_reset_reset_bridge_in_reset.reset
		.master_jtag_master_address                                               (master_jtag_master_address),                                         //                                                 master_jtag_master.address
		.master_jtag_master_waitrequest                                           (master_jtag_master_waitrequest),                                     //                                                                   .waitrequest
		.master_jtag_master_byteenable                                            (master_jtag_master_byteenable),                                      //                                                                   .byteenable
		.master_jtag_master_read                                                  (master_jtag_master_read),                                            //                                                                   .read
		.master_jtag_master_readdata                                              (master_jtag_master_readdata),                                        //                                                                   .readdata
		.master_jtag_master_readdatavalid                                         (master_jtag_master_readdatavalid),                                   //                                                                   .readdatavalid
		.master_jtag_master_write                                                 (master_jtag_master_write),                                           //                                                                   .write
		.master_jtag_master_writedata                                             (master_jtag_master_writedata),                                       //                                                                   .writedata
		.a_4_quadrant_chopper_0_avalon_slave_0_address                            (mm_interconnect_0_a_4_quadrant_chopper_0_avalon_slave_0_address),    //                              a_4_quadrant_chopper_0_avalon_slave_0.address
		.a_4_quadrant_chopper_0_avalon_slave_0_write                              (mm_interconnect_0_a_4_quadrant_chopper_0_avalon_slave_0_write),      //                                                                   .write
		.a_4_quadrant_chopper_0_avalon_slave_0_read                               (mm_interconnect_0_a_4_quadrant_chopper_0_avalon_slave_0_read),       //                                                                   .read
		.a_4_quadrant_chopper_0_avalon_slave_0_readdata                           (mm_interconnect_0_a_4_quadrant_chopper_0_avalon_slave_0_readdata),   //                                                                   .readdata
		.a_4_quadrant_chopper_0_avalon_slave_0_writedata                          (mm_interconnect_0_a_4_quadrant_chopper_0_avalon_slave_0_writedata),  //                                                                   .writedata
		.a_4_quadrant_chopper_0_avalon_slave_0_byteenable                         (mm_interconnect_0_a_4_quadrant_chopper_0_avalon_slave_0_byteenable), //                                                                   .byteenable
		.sysid_control_slave_address                                              (mm_interconnect_0_sysid_control_slave_address),                      //                                                sysid_control_slave.address
		.sysid_control_slave_readdata                                             (mm_interconnect_0_sysid_control_slave_readdata)                      //                                                                   .readdata
	);

	core_irq_mapper irq_mapper (
		.clk           (),                          //       clk.clk
		.reset         (),                          // clk_reset.reset
		.receiver0_irq (~irq_mapper_receiver0_irq), // receiver0.irq
		.sender_irq    (hps_system_f2h_irq0_irq)    //    sender.irq
	);

	core_irq_mapper_001 irq_mapper_001 (
		.clk        (),                        //       clk.clk
		.reset      (),                        // clk_reset.reset
		.sender_irq (hps_system_f2h_irq1_irq)  //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (pll_0_outclk0_clk),              //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~hps_system_h2f_reset_reset),        // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
