-- core.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity core is
	port (
		clk_clk                         : in    std_logic                     := '0';             --    clk.clk
		hps_io_hps_io_emac1_inst_TX_CLK : out   std_logic;                                        -- hps_io.hps_io_emac1_inst_TX_CLK
		hps_io_hps_io_emac1_inst_TXD0   : out   std_logic;                                        --       .hps_io_emac1_inst_TXD0
		hps_io_hps_io_emac1_inst_TXD1   : out   std_logic;                                        --       .hps_io_emac1_inst_TXD1
		hps_io_hps_io_emac1_inst_TXD2   : out   std_logic;                                        --       .hps_io_emac1_inst_TXD2
		hps_io_hps_io_emac1_inst_TXD3   : out   std_logic;                                        --       .hps_io_emac1_inst_TXD3
		hps_io_hps_io_emac1_inst_RXD0   : in    std_logic                     := '0';             --       .hps_io_emac1_inst_RXD0
		hps_io_hps_io_emac1_inst_MDIO   : inout std_logic                     := '0';             --       .hps_io_emac1_inst_MDIO
		hps_io_hps_io_emac1_inst_MDC    : out   std_logic;                                        --       .hps_io_emac1_inst_MDC
		hps_io_hps_io_emac1_inst_RX_CTL : in    std_logic                     := '0';             --       .hps_io_emac1_inst_RX_CTL
		hps_io_hps_io_emac1_inst_TX_CTL : out   std_logic;                                        --       .hps_io_emac1_inst_TX_CTL
		hps_io_hps_io_emac1_inst_RX_CLK : in    std_logic                     := '0';             --       .hps_io_emac1_inst_RX_CLK
		hps_io_hps_io_emac1_inst_RXD1   : in    std_logic                     := '0';             --       .hps_io_emac1_inst_RXD1
		hps_io_hps_io_emac1_inst_RXD2   : in    std_logic                     := '0';             --       .hps_io_emac1_inst_RXD2
		hps_io_hps_io_emac1_inst_RXD3   : in    std_logic                     := '0';             --       .hps_io_emac1_inst_RXD3
		hps_io_hps_io_sdio_inst_CMD     : inout std_logic                     := '0';             --       .hps_io_sdio_inst_CMD
		hps_io_hps_io_sdio_inst_D0      : inout std_logic                     := '0';             --       .hps_io_sdio_inst_D0
		hps_io_hps_io_sdio_inst_D1      : inout std_logic                     := '0';             --       .hps_io_sdio_inst_D1
		hps_io_hps_io_sdio_inst_CLK     : out   std_logic;                                        --       .hps_io_sdio_inst_CLK
		hps_io_hps_io_sdio_inst_D2      : inout std_logic                     := '0';             --       .hps_io_sdio_inst_D2
		hps_io_hps_io_sdio_inst_D3      : inout std_logic                     := '0';             --       .hps_io_sdio_inst_D3
		hps_io_hps_io_uart0_inst_RX     : in    std_logic                     := '0';             --       .hps_io_uart0_inst_RX
		hps_io_hps_io_uart0_inst_TX     : out   std_logic;                                        --       .hps_io_uart0_inst_TX
		hps_io_hps_io_i2c0_inst_SDA     : inout std_logic                     := '0';             --       .hps_io_i2c0_inst_SDA
		hps_io_hps_io_i2c0_inst_SCL     : inout std_logic                     := '0';             --       .hps_io_i2c0_inst_SCL
		hps_io_hps_io_i2c1_inst_SDA     : inout std_logic                     := '0';             --       .hps_io_i2c1_inst_SDA
		hps_io_hps_io_i2c1_inst_SCL     : inout std_logic                     := '0';             --       .hps_io_i2c1_inst_SCL
		memory_mem_a                    : out   std_logic_vector(14 downto 0);                    -- memory.mem_a
		memory_mem_ba                   : out   std_logic_vector(2 downto 0);                     --       .mem_ba
		memory_mem_ck                   : out   std_logic;                                        --       .mem_ck
		memory_mem_ck_n                 : out   std_logic;                                        --       .mem_ck_n
		memory_mem_cke                  : out   std_logic;                                        --       .mem_cke
		memory_mem_cs_n                 : out   std_logic;                                        --       .mem_cs_n
		memory_mem_ras_n                : out   std_logic;                                        --       .mem_ras_n
		memory_mem_cas_n                : out   std_logic;                                        --       .mem_cas_n
		memory_mem_we_n                 : out   std_logic;                                        --       .mem_we_n
		memory_mem_reset_n              : out   std_logic;                                        --       .mem_reset_n
		memory_mem_dq                   : inout std_logic_vector(31 downto 0) := (others => '0'); --       .mem_dq
		memory_mem_dqs                  : inout std_logic_vector(3 downto 0)  := (others => '0'); --       .mem_dqs
		memory_mem_dqs_n                : inout std_logic_vector(3 downto 0)  := (others => '0'); --       .mem_dqs_n
		memory_mem_odt                  : out   std_logic;                                        --       .mem_odt
		memory_mem_dm                   : out   std_logic_vector(3 downto 0);                     --       .mem_dm
		memory_oct_rzqin                : in    std_logic                     := '0';             --       .oct_rzqin
		pwm_a_pwm                       : out   std_logic;                                        --    pwm.a_pwm
		pwm_b_pwm                       : out   std_logic;                                        --       .b_pwm
		pwm_secure                      : in    std_logic                     := '0';             --       .secure
		reset_reset_n                   : in    std_logic                     := '0'              --  reset.reset_n
	);
end entity core;

architecture rtl of core is
	component hacheur_top is
		port (
			rsi_reset      : in  std_logic                     := 'X';             -- reset
			avs_address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			avs_byteenable : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable
			avs_read       : in  std_logic                     := 'X';             -- read
			avs_readdata   : out std_logic_vector(15 downto 0);                    -- readdata
			avs_write      : in  std_logic                     := 'X';             -- write
			avs_writedata  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			ins_end_cycle  : out std_logic;                                        -- irq_n
			csi_clock      : in  std_logic                     := 'X';             -- clk
			A              : out std_logic;                                        -- a_pwm
			B              : out std_logic;                                        -- b_pwm
			secure         : in  std_logic                     := 'X'              -- secure
		);
	end component hacheur_top;

	component core_hps_system is
		generic (
			F2S_Width : integer := 2;
			S2F_Width : integer := 2
		);
		port (
			h2f_mpu_eventi           : in    std_logic                     := 'X';             -- eventi
			h2f_mpu_evento           : out   std_logic;                                        -- evento
			h2f_mpu_standbywfe       : out   std_logic_vector(1 downto 0);                     -- standbywfe
			h2f_mpu_standbywfi       : out   std_logic_vector(1 downto 0);                     -- standbywfi
			mem_a                    : out   std_logic_vector(14 downto 0);                    -- mem_a
			mem_ba                   : out   std_logic_vector(2 downto 0);                     -- mem_ba
			mem_ck                   : out   std_logic;                                        -- mem_ck
			mem_ck_n                 : out   std_logic;                                        -- mem_ck_n
			mem_cke                  : out   std_logic;                                        -- mem_cke
			mem_cs_n                 : out   std_logic;                                        -- mem_cs_n
			mem_ras_n                : out   std_logic;                                        -- mem_ras_n
			mem_cas_n                : out   std_logic;                                        -- mem_cas_n
			mem_we_n                 : out   std_logic;                                        -- mem_we_n
			mem_reset_n              : out   std_logic;                                        -- mem_reset_n
			mem_dq                   : inout std_logic_vector(31 downto 0) := (others => 'X'); -- mem_dq
			mem_dqs                  : inout std_logic_vector(3 downto 0)  := (others => 'X'); -- mem_dqs
			mem_dqs_n                : inout std_logic_vector(3 downto 0)  := (others => 'X'); -- mem_dqs_n
			mem_odt                  : out   std_logic;                                        -- mem_odt
			mem_dm                   : out   std_logic_vector(3 downto 0);                     -- mem_dm
			oct_rzqin                : in    std_logic                     := 'X';             -- oct_rzqin
			hps_io_emac1_inst_TX_CLK : out   std_logic;                                        -- hps_io_emac1_inst_TX_CLK
			hps_io_emac1_inst_TXD0   : out   std_logic;                                        -- hps_io_emac1_inst_TXD0
			hps_io_emac1_inst_TXD1   : out   std_logic;                                        -- hps_io_emac1_inst_TXD1
			hps_io_emac1_inst_TXD2   : out   std_logic;                                        -- hps_io_emac1_inst_TXD2
			hps_io_emac1_inst_TXD3   : out   std_logic;                                        -- hps_io_emac1_inst_TXD3
			hps_io_emac1_inst_RXD0   : in    std_logic                     := 'X';             -- hps_io_emac1_inst_RXD0
			hps_io_emac1_inst_MDIO   : inout std_logic                     := 'X';             -- hps_io_emac1_inst_MDIO
			hps_io_emac1_inst_MDC    : out   std_logic;                                        -- hps_io_emac1_inst_MDC
			hps_io_emac1_inst_RX_CTL : in    std_logic                     := 'X';             -- hps_io_emac1_inst_RX_CTL
			hps_io_emac1_inst_TX_CTL : out   std_logic;                                        -- hps_io_emac1_inst_TX_CTL
			hps_io_emac1_inst_RX_CLK : in    std_logic                     := 'X';             -- hps_io_emac1_inst_RX_CLK
			hps_io_emac1_inst_RXD1   : in    std_logic                     := 'X';             -- hps_io_emac1_inst_RXD1
			hps_io_emac1_inst_RXD2   : in    std_logic                     := 'X';             -- hps_io_emac1_inst_RXD2
			hps_io_emac1_inst_RXD3   : in    std_logic                     := 'X';             -- hps_io_emac1_inst_RXD3
			hps_io_sdio_inst_CMD     : inout std_logic                     := 'X';             -- hps_io_sdio_inst_CMD
			hps_io_sdio_inst_D0      : inout std_logic                     := 'X';             -- hps_io_sdio_inst_D0
			hps_io_sdio_inst_D1      : inout std_logic                     := 'X';             -- hps_io_sdio_inst_D1
			hps_io_sdio_inst_CLK     : out   std_logic;                                        -- hps_io_sdio_inst_CLK
			hps_io_sdio_inst_D2      : inout std_logic                     := 'X';             -- hps_io_sdio_inst_D2
			hps_io_sdio_inst_D3      : inout std_logic                     := 'X';             -- hps_io_sdio_inst_D3
			hps_io_uart0_inst_RX     : in    std_logic                     := 'X';             -- hps_io_uart0_inst_RX
			hps_io_uart0_inst_TX     : out   std_logic;                                        -- hps_io_uart0_inst_TX
			hps_io_i2c0_inst_SDA     : inout std_logic                     := 'X';             -- hps_io_i2c0_inst_SDA
			hps_io_i2c0_inst_SCL     : inout std_logic                     := 'X';             -- hps_io_i2c0_inst_SCL
			hps_io_i2c1_inst_SDA     : inout std_logic                     := 'X';             -- hps_io_i2c1_inst_SDA
			hps_io_i2c1_inst_SCL     : inout std_logic                     := 'X';             -- hps_io_i2c1_inst_SCL
			h2f_rst_n                : out   std_logic;                                        -- reset_n
			f2h_sdram0_clk           : in    std_logic                     := 'X';             -- clk
			f2h_sdram0_ARADDR        : in    std_logic_vector(31 downto 0) := (others => 'X'); -- araddr
			f2h_sdram0_ARLEN         : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- arlen
			f2h_sdram0_ARID          : in    std_logic_vector(7 downto 0)  := (others => 'X'); -- arid
			f2h_sdram0_ARSIZE        : in    std_logic_vector(2 downto 0)  := (others => 'X'); -- arsize
			f2h_sdram0_ARBURST       : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- arburst
			f2h_sdram0_ARLOCK        : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- arlock
			f2h_sdram0_ARPROT        : in    std_logic_vector(2 downto 0)  := (others => 'X'); -- arprot
			f2h_sdram0_ARVALID       : in    std_logic                     := 'X';             -- arvalid
			f2h_sdram0_ARCACHE       : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- arcache
			f2h_sdram0_AWADDR        : in    std_logic_vector(31 downto 0) := (others => 'X'); -- awaddr
			f2h_sdram0_AWLEN         : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- awlen
			f2h_sdram0_AWID          : in    std_logic_vector(7 downto 0)  := (others => 'X'); -- awid
			f2h_sdram0_AWSIZE        : in    std_logic_vector(2 downto 0)  := (others => 'X'); -- awsize
			f2h_sdram0_AWBURST       : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- awburst
			f2h_sdram0_AWLOCK        : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- awlock
			f2h_sdram0_AWPROT        : in    std_logic_vector(2 downto 0)  := (others => 'X'); -- awprot
			f2h_sdram0_AWVALID       : in    std_logic                     := 'X';             -- awvalid
			f2h_sdram0_AWCACHE       : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- awcache
			f2h_sdram0_BRESP         : out   std_logic_vector(1 downto 0);                     -- bresp
			f2h_sdram0_BID           : out   std_logic_vector(7 downto 0);                     -- bid
			f2h_sdram0_BVALID        : out   std_logic;                                        -- bvalid
			f2h_sdram0_BREADY        : in    std_logic                     := 'X';             -- bready
			f2h_sdram0_ARREADY       : out   std_logic;                                        -- arready
			f2h_sdram0_AWREADY       : out   std_logic;                                        -- awready
			f2h_sdram0_RREADY        : in    std_logic                     := 'X';             -- rready
			f2h_sdram0_RDATA         : out   std_logic_vector(63 downto 0);                    -- rdata
			f2h_sdram0_RRESP         : out   std_logic_vector(1 downto 0);                     -- rresp
			f2h_sdram0_RLAST         : out   std_logic;                                        -- rlast
			f2h_sdram0_RID           : out   std_logic_vector(7 downto 0);                     -- rid
			f2h_sdram0_RVALID        : out   std_logic;                                        -- rvalid
			f2h_sdram0_WLAST         : in    std_logic                     := 'X';             -- wlast
			f2h_sdram0_WVALID        : in    std_logic                     := 'X';             -- wvalid
			f2h_sdram0_WDATA         : in    std_logic_vector(63 downto 0) := (others => 'X'); -- wdata
			f2h_sdram0_WSTRB         : in    std_logic_vector(7 downto 0)  := (others => 'X'); -- wstrb
			f2h_sdram0_WREADY        : out   std_logic;                                        -- wready
			f2h_sdram0_WID           : in    std_logic_vector(7 downto 0)  := (others => 'X'); -- wid
			h2f_axi_clk              : in    std_logic                     := 'X';             -- clk
			h2f_AWID                 : out   std_logic_vector(11 downto 0);                    -- awid
			h2f_AWADDR               : out   std_logic_vector(29 downto 0);                    -- awaddr
			h2f_AWLEN                : out   std_logic_vector(3 downto 0);                     -- awlen
			h2f_AWSIZE               : out   std_logic_vector(2 downto 0);                     -- awsize
			h2f_AWBURST              : out   std_logic_vector(1 downto 0);                     -- awburst
			h2f_AWLOCK               : out   std_logic_vector(1 downto 0);                     -- awlock
			h2f_AWCACHE              : out   std_logic_vector(3 downto 0);                     -- awcache
			h2f_AWPROT               : out   std_logic_vector(2 downto 0);                     -- awprot
			h2f_AWVALID              : out   std_logic;                                        -- awvalid
			h2f_AWREADY              : in    std_logic                     := 'X';             -- awready
			h2f_WID                  : out   std_logic_vector(11 downto 0);                    -- wid
			h2f_WDATA                : out   std_logic_vector(63 downto 0);                    -- wdata
			h2f_WSTRB                : out   std_logic_vector(7 downto 0);                     -- wstrb
			h2f_WLAST                : out   std_logic;                                        -- wlast
			h2f_WVALID               : out   std_logic;                                        -- wvalid
			h2f_WREADY               : in    std_logic                     := 'X';             -- wready
			h2f_BID                  : in    std_logic_vector(11 downto 0) := (others => 'X'); -- bid
			h2f_BRESP                : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- bresp
			h2f_BVALID               : in    std_logic                     := 'X';             -- bvalid
			h2f_BREADY               : out   std_logic;                                        -- bready
			h2f_ARID                 : out   std_logic_vector(11 downto 0);                    -- arid
			h2f_ARADDR               : out   std_logic_vector(29 downto 0);                    -- araddr
			h2f_ARLEN                : out   std_logic_vector(3 downto 0);                     -- arlen
			h2f_ARSIZE               : out   std_logic_vector(2 downto 0);                     -- arsize
			h2f_ARBURST              : out   std_logic_vector(1 downto 0);                     -- arburst
			h2f_ARLOCK               : out   std_logic_vector(1 downto 0);                     -- arlock
			h2f_ARCACHE              : out   std_logic_vector(3 downto 0);                     -- arcache
			h2f_ARPROT               : out   std_logic_vector(2 downto 0);                     -- arprot
			h2f_ARVALID              : out   std_logic;                                        -- arvalid
			h2f_ARREADY              : in    std_logic                     := 'X';             -- arready
			h2f_RID                  : in    std_logic_vector(11 downto 0) := (others => 'X'); -- rid
			h2f_RDATA                : in    std_logic_vector(63 downto 0) := (others => 'X'); -- rdata
			h2f_RRESP                : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- rresp
			h2f_RLAST                : in    std_logic                     := 'X';             -- rlast
			h2f_RVALID               : in    std_logic                     := 'X';             -- rvalid
			h2f_RREADY               : out   std_logic;                                        -- rready
			f2h_axi_clk              : in    std_logic                     := 'X';             -- clk
			f2h_AWID                 : in    std_logic_vector(7 downto 0)  := (others => 'X'); -- awid
			f2h_AWADDR               : in    std_logic_vector(31 downto 0) := (others => 'X'); -- awaddr
			f2h_AWLEN                : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- awlen
			f2h_AWSIZE               : in    std_logic_vector(2 downto 0)  := (others => 'X'); -- awsize
			f2h_AWBURST              : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- awburst
			f2h_AWLOCK               : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- awlock
			f2h_AWCACHE              : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- awcache
			f2h_AWPROT               : in    std_logic_vector(2 downto 0)  := (others => 'X'); -- awprot
			f2h_AWVALID              : in    std_logic                     := 'X';             -- awvalid
			f2h_AWREADY              : out   std_logic;                                        -- awready
			f2h_AWUSER               : in    std_logic_vector(4 downto 0)  := (others => 'X'); -- awuser
			f2h_WID                  : in    std_logic_vector(7 downto 0)  := (others => 'X'); -- wid
			f2h_WDATA                : in    std_logic_vector(63 downto 0) := (others => 'X'); -- wdata
			f2h_WSTRB                : in    std_logic_vector(7 downto 0)  := (others => 'X'); -- wstrb
			f2h_WLAST                : in    std_logic                     := 'X';             -- wlast
			f2h_WVALID               : in    std_logic                     := 'X';             -- wvalid
			f2h_WREADY               : out   std_logic;                                        -- wready
			f2h_BID                  : out   std_logic_vector(7 downto 0);                     -- bid
			f2h_BRESP                : out   std_logic_vector(1 downto 0);                     -- bresp
			f2h_BVALID               : out   std_logic;                                        -- bvalid
			f2h_BREADY               : in    std_logic                     := 'X';             -- bready
			f2h_ARID                 : in    std_logic_vector(7 downto 0)  := (others => 'X'); -- arid
			f2h_ARADDR               : in    std_logic_vector(31 downto 0) := (others => 'X'); -- araddr
			f2h_ARLEN                : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- arlen
			f2h_ARSIZE               : in    std_logic_vector(2 downto 0)  := (others => 'X'); -- arsize
			f2h_ARBURST              : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- arburst
			f2h_ARLOCK               : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- arlock
			f2h_ARCACHE              : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- arcache
			f2h_ARPROT               : in    std_logic_vector(2 downto 0)  := (others => 'X'); -- arprot
			f2h_ARVALID              : in    std_logic                     := 'X';             -- arvalid
			f2h_ARREADY              : out   std_logic;                                        -- arready
			f2h_ARUSER               : in    std_logic_vector(4 downto 0)  := (others => 'X'); -- aruser
			f2h_RID                  : out   std_logic_vector(7 downto 0);                     -- rid
			f2h_RDATA                : out   std_logic_vector(63 downto 0);                    -- rdata
			f2h_RRESP                : out   std_logic_vector(1 downto 0);                     -- rresp
			f2h_RLAST                : out   std_logic;                                        -- rlast
			f2h_RVALID               : out   std_logic;                                        -- rvalid
			f2h_RREADY               : in    std_logic                     := 'X';             -- rready
			h2f_lw_axi_clk           : in    std_logic                     := 'X';             -- clk
			h2f_lw_AWID              : out   std_logic_vector(11 downto 0);                    -- awid
			h2f_lw_AWADDR            : out   std_logic_vector(20 downto 0);                    -- awaddr
			h2f_lw_AWLEN             : out   std_logic_vector(3 downto 0);                     -- awlen
			h2f_lw_AWSIZE            : out   std_logic_vector(2 downto 0);                     -- awsize
			h2f_lw_AWBURST           : out   std_logic_vector(1 downto 0);                     -- awburst
			h2f_lw_AWLOCK            : out   std_logic_vector(1 downto 0);                     -- awlock
			h2f_lw_AWCACHE           : out   std_logic_vector(3 downto 0);                     -- awcache
			h2f_lw_AWPROT            : out   std_logic_vector(2 downto 0);                     -- awprot
			h2f_lw_AWVALID           : out   std_logic;                                        -- awvalid
			h2f_lw_AWREADY           : in    std_logic                     := 'X';             -- awready
			h2f_lw_WID               : out   std_logic_vector(11 downto 0);                    -- wid
			h2f_lw_WDATA             : out   std_logic_vector(31 downto 0);                    -- wdata
			h2f_lw_WSTRB             : out   std_logic_vector(3 downto 0);                     -- wstrb
			h2f_lw_WLAST             : out   std_logic;                                        -- wlast
			h2f_lw_WVALID            : out   std_logic;                                        -- wvalid
			h2f_lw_WREADY            : in    std_logic                     := 'X';             -- wready
			h2f_lw_BID               : in    std_logic_vector(11 downto 0) := (others => 'X'); -- bid
			h2f_lw_BRESP             : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- bresp
			h2f_lw_BVALID            : in    std_logic                     := 'X';             -- bvalid
			h2f_lw_BREADY            : out   std_logic;                                        -- bready
			h2f_lw_ARID              : out   std_logic_vector(11 downto 0);                    -- arid
			h2f_lw_ARADDR            : out   std_logic_vector(20 downto 0);                    -- araddr
			h2f_lw_ARLEN             : out   std_logic_vector(3 downto 0);                     -- arlen
			h2f_lw_ARSIZE            : out   std_logic_vector(2 downto 0);                     -- arsize
			h2f_lw_ARBURST           : out   std_logic_vector(1 downto 0);                     -- arburst
			h2f_lw_ARLOCK            : out   std_logic_vector(1 downto 0);                     -- arlock
			h2f_lw_ARCACHE           : out   std_logic_vector(3 downto 0);                     -- arcache
			h2f_lw_ARPROT            : out   std_logic_vector(2 downto 0);                     -- arprot
			h2f_lw_ARVALID           : out   std_logic;                                        -- arvalid
			h2f_lw_ARREADY           : in    std_logic                     := 'X';             -- arready
			h2f_lw_RID               : in    std_logic_vector(11 downto 0) := (others => 'X'); -- rid
			h2f_lw_RDATA             : in    std_logic_vector(31 downto 0) := (others => 'X'); -- rdata
			h2f_lw_RRESP             : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- rresp
			h2f_lw_RLAST             : in    std_logic                     := 'X';             -- rlast
			h2f_lw_RVALID            : in    std_logic                     := 'X';             -- rvalid
			h2f_lw_RREADY            : out   std_logic;                                        -- rready
			f2h_irq_p0               : in    std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			f2h_irq_p1               : in    std_logic_vector(31 downto 0) := (others => 'X')  -- irq
		);
	end component core_hps_system;

	component core_master_jtag is
		generic (
			USE_PLI     : integer := 0;
			PLI_PORT    : integer := 50000;
			FIFO_DEPTHS : integer := 2
		);
		port (
			clk_clk              : in  std_logic                     := 'X';             -- clk
			clk_reset_reset      : in  std_logic                     := 'X';             -- reset
			master_address       : out std_logic_vector(31 downto 0);                    -- address
			master_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			master_read          : out std_logic;                                        -- read
			master_write         : out std_logic;                                        -- write
			master_writedata     : out std_logic_vector(31 downto 0);                    -- writedata
			master_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			master_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			master_byteenable    : out std_logic_vector(3 downto 0);                     -- byteenable
			master_reset_reset   : out std_logic                                         -- reset
		);
	end component core_master_jtag;

	component core_sysid is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component core_sysid;

	component core_mm_interconnect_0 is
		port (
			hps_system_h2f_lw_axi_master_awid                                        : in  std_logic_vector(11 downto 0) := (others => 'X'); -- awid
			hps_system_h2f_lw_axi_master_awaddr                                      : in  std_logic_vector(20 downto 0) := (others => 'X'); -- awaddr
			hps_system_h2f_lw_axi_master_awlen                                       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- awlen
			hps_system_h2f_lw_axi_master_awsize                                      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- awsize
			hps_system_h2f_lw_axi_master_awburst                                     : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- awburst
			hps_system_h2f_lw_axi_master_awlock                                      : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- awlock
			hps_system_h2f_lw_axi_master_awcache                                     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- awcache
			hps_system_h2f_lw_axi_master_awprot                                      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- awprot
			hps_system_h2f_lw_axi_master_awvalid                                     : in  std_logic                     := 'X';             -- awvalid
			hps_system_h2f_lw_axi_master_awready                                     : out std_logic;                                        -- awready
			hps_system_h2f_lw_axi_master_wid                                         : in  std_logic_vector(11 downto 0) := (others => 'X'); -- wid
			hps_system_h2f_lw_axi_master_wdata                                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- wdata
			hps_system_h2f_lw_axi_master_wstrb                                       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- wstrb
			hps_system_h2f_lw_axi_master_wlast                                       : in  std_logic                     := 'X';             -- wlast
			hps_system_h2f_lw_axi_master_wvalid                                      : in  std_logic                     := 'X';             -- wvalid
			hps_system_h2f_lw_axi_master_wready                                      : out std_logic;                                        -- wready
			hps_system_h2f_lw_axi_master_bid                                         : out std_logic_vector(11 downto 0);                    -- bid
			hps_system_h2f_lw_axi_master_bresp                                       : out std_logic_vector(1 downto 0);                     -- bresp
			hps_system_h2f_lw_axi_master_bvalid                                      : out std_logic;                                        -- bvalid
			hps_system_h2f_lw_axi_master_bready                                      : in  std_logic                     := 'X';             -- bready
			hps_system_h2f_lw_axi_master_arid                                        : in  std_logic_vector(11 downto 0) := (others => 'X'); -- arid
			hps_system_h2f_lw_axi_master_araddr                                      : in  std_logic_vector(20 downto 0) := (others => 'X'); -- araddr
			hps_system_h2f_lw_axi_master_arlen                                       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- arlen
			hps_system_h2f_lw_axi_master_arsize                                      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- arsize
			hps_system_h2f_lw_axi_master_arburst                                     : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- arburst
			hps_system_h2f_lw_axi_master_arlock                                      : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- arlock
			hps_system_h2f_lw_axi_master_arcache                                     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- arcache
			hps_system_h2f_lw_axi_master_arprot                                      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- arprot
			hps_system_h2f_lw_axi_master_arvalid                                     : in  std_logic                     := 'X';             -- arvalid
			hps_system_h2f_lw_axi_master_arready                                     : out std_logic;                                        -- arready
			hps_system_h2f_lw_axi_master_rid                                         : out std_logic_vector(11 downto 0);                    -- rid
			hps_system_h2f_lw_axi_master_rdata                                       : out std_logic_vector(31 downto 0);                    -- rdata
			hps_system_h2f_lw_axi_master_rresp                                       : out std_logic_vector(1 downto 0);                     -- rresp
			hps_system_h2f_lw_axi_master_rlast                                       : out std_logic;                                        -- rlast
			hps_system_h2f_lw_axi_master_rvalid                                      : out std_logic;                                        -- rvalid
			hps_system_h2f_lw_axi_master_rready                                      : in  std_logic                     := 'X';             -- rready
			clk_0_clk_clk                                                            : in  std_logic                     := 'X';             -- clk
			a_4_quadrant_chopper_0_clock_reset_reset_bridge_in_reset_reset           : in  std_logic                     := 'X';             -- reset
			hps_system_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			master_jtag_clk_reset_reset_bridge_in_reset_reset                        : in  std_logic                     := 'X';             -- reset
			master_jtag_master_address                                               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			master_jtag_master_waitrequest                                           : out std_logic;                                        -- waitrequest
			master_jtag_master_byteenable                                            : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			master_jtag_master_read                                                  : in  std_logic                     := 'X';             -- read
			master_jtag_master_readdata                                              : out std_logic_vector(31 downto 0);                    -- readdata
			master_jtag_master_readdatavalid                                         : out std_logic;                                        -- readdatavalid
			master_jtag_master_write                                                 : in  std_logic                     := 'X';             -- write
			master_jtag_master_writedata                                             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			a_4_quadrant_chopper_0_avalon_slave_0_address                            : out std_logic_vector(1 downto 0);                     -- address
			a_4_quadrant_chopper_0_avalon_slave_0_write                              : out std_logic;                                        -- write
			a_4_quadrant_chopper_0_avalon_slave_0_read                               : out std_logic;                                        -- read
			a_4_quadrant_chopper_0_avalon_slave_0_readdata                           : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			a_4_quadrant_chopper_0_avalon_slave_0_writedata                          : out std_logic_vector(15 downto 0);                    -- writedata
			a_4_quadrant_chopper_0_avalon_slave_0_byteenable                         : out std_logic_vector(1 downto 0);                     -- byteenable
			sysid_control_slave_address                                              : out std_logic_vector(0 downto 0);                     -- address
			sysid_control_slave_readdata                                             : in  std_logic_vector(31 downto 0) := (others => 'X')  -- readdata
		);
	end component core_mm_interconnect_0;

	component core_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component core_irq_mapper;

	component core_irq_mapper_001 is
		port (
			clk        : in  std_logic                     := 'X'; -- clk
			reset      : in  std_logic                     := 'X'; -- reset
			sender_irq : out std_logic_vector(31 downto 0)         -- irq
		);
	end component core_irq_mapper_001;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component altera_reset_controller;

	signal hps_system_h2f_lw_axi_master_awburst                               : std_logic_vector(1 downto 0);  -- hps_system:h2f_lw_AWBURST -> mm_interconnect_0:hps_system_h2f_lw_axi_master_awburst
	signal hps_system_h2f_lw_axi_master_arlen                                 : std_logic_vector(3 downto 0);  -- hps_system:h2f_lw_ARLEN -> mm_interconnect_0:hps_system_h2f_lw_axi_master_arlen
	signal hps_system_h2f_lw_axi_master_wstrb                                 : std_logic_vector(3 downto 0);  -- hps_system:h2f_lw_WSTRB -> mm_interconnect_0:hps_system_h2f_lw_axi_master_wstrb
	signal hps_system_h2f_lw_axi_master_wready                                : std_logic;                     -- mm_interconnect_0:hps_system_h2f_lw_axi_master_wready -> hps_system:h2f_lw_WREADY
	signal hps_system_h2f_lw_axi_master_rid                                   : std_logic_vector(11 downto 0); -- mm_interconnect_0:hps_system_h2f_lw_axi_master_rid -> hps_system:h2f_lw_RID
	signal hps_system_h2f_lw_axi_master_rready                                : std_logic;                     -- hps_system:h2f_lw_RREADY -> mm_interconnect_0:hps_system_h2f_lw_axi_master_rready
	signal hps_system_h2f_lw_axi_master_awlen                                 : std_logic_vector(3 downto 0);  -- hps_system:h2f_lw_AWLEN -> mm_interconnect_0:hps_system_h2f_lw_axi_master_awlen
	signal hps_system_h2f_lw_axi_master_wid                                   : std_logic_vector(11 downto 0); -- hps_system:h2f_lw_WID -> mm_interconnect_0:hps_system_h2f_lw_axi_master_wid
	signal hps_system_h2f_lw_axi_master_arcache                               : std_logic_vector(3 downto 0);  -- hps_system:h2f_lw_ARCACHE -> mm_interconnect_0:hps_system_h2f_lw_axi_master_arcache
	signal hps_system_h2f_lw_axi_master_wvalid                                : std_logic;                     -- hps_system:h2f_lw_WVALID -> mm_interconnect_0:hps_system_h2f_lw_axi_master_wvalid
	signal hps_system_h2f_lw_axi_master_araddr                                : std_logic_vector(20 downto 0); -- hps_system:h2f_lw_ARADDR -> mm_interconnect_0:hps_system_h2f_lw_axi_master_araddr
	signal hps_system_h2f_lw_axi_master_arprot                                : std_logic_vector(2 downto 0);  -- hps_system:h2f_lw_ARPROT -> mm_interconnect_0:hps_system_h2f_lw_axi_master_arprot
	signal hps_system_h2f_lw_axi_master_awprot                                : std_logic_vector(2 downto 0);  -- hps_system:h2f_lw_AWPROT -> mm_interconnect_0:hps_system_h2f_lw_axi_master_awprot
	signal hps_system_h2f_lw_axi_master_wdata                                 : std_logic_vector(31 downto 0); -- hps_system:h2f_lw_WDATA -> mm_interconnect_0:hps_system_h2f_lw_axi_master_wdata
	signal hps_system_h2f_lw_axi_master_arvalid                               : std_logic;                     -- hps_system:h2f_lw_ARVALID -> mm_interconnect_0:hps_system_h2f_lw_axi_master_arvalid
	signal hps_system_h2f_lw_axi_master_awcache                               : std_logic_vector(3 downto 0);  -- hps_system:h2f_lw_AWCACHE -> mm_interconnect_0:hps_system_h2f_lw_axi_master_awcache
	signal hps_system_h2f_lw_axi_master_arid                                  : std_logic_vector(11 downto 0); -- hps_system:h2f_lw_ARID -> mm_interconnect_0:hps_system_h2f_lw_axi_master_arid
	signal hps_system_h2f_lw_axi_master_arlock                                : std_logic_vector(1 downto 0);  -- hps_system:h2f_lw_ARLOCK -> mm_interconnect_0:hps_system_h2f_lw_axi_master_arlock
	signal hps_system_h2f_lw_axi_master_awlock                                : std_logic_vector(1 downto 0);  -- hps_system:h2f_lw_AWLOCK -> mm_interconnect_0:hps_system_h2f_lw_axi_master_awlock
	signal hps_system_h2f_lw_axi_master_awaddr                                : std_logic_vector(20 downto 0); -- hps_system:h2f_lw_AWADDR -> mm_interconnect_0:hps_system_h2f_lw_axi_master_awaddr
	signal hps_system_h2f_lw_axi_master_bresp                                 : std_logic_vector(1 downto 0);  -- mm_interconnect_0:hps_system_h2f_lw_axi_master_bresp -> hps_system:h2f_lw_BRESP
	signal hps_system_h2f_lw_axi_master_arready                               : std_logic;                     -- mm_interconnect_0:hps_system_h2f_lw_axi_master_arready -> hps_system:h2f_lw_ARREADY
	signal hps_system_h2f_lw_axi_master_rdata                                 : std_logic_vector(31 downto 0); -- mm_interconnect_0:hps_system_h2f_lw_axi_master_rdata -> hps_system:h2f_lw_RDATA
	signal hps_system_h2f_lw_axi_master_awready                               : std_logic;                     -- mm_interconnect_0:hps_system_h2f_lw_axi_master_awready -> hps_system:h2f_lw_AWREADY
	signal hps_system_h2f_lw_axi_master_arburst                               : std_logic_vector(1 downto 0);  -- hps_system:h2f_lw_ARBURST -> mm_interconnect_0:hps_system_h2f_lw_axi_master_arburst
	signal hps_system_h2f_lw_axi_master_arsize                                : std_logic_vector(2 downto 0);  -- hps_system:h2f_lw_ARSIZE -> mm_interconnect_0:hps_system_h2f_lw_axi_master_arsize
	signal hps_system_h2f_lw_axi_master_bready                                : std_logic;                     -- hps_system:h2f_lw_BREADY -> mm_interconnect_0:hps_system_h2f_lw_axi_master_bready
	signal hps_system_h2f_lw_axi_master_rlast                                 : std_logic;                     -- mm_interconnect_0:hps_system_h2f_lw_axi_master_rlast -> hps_system:h2f_lw_RLAST
	signal hps_system_h2f_lw_axi_master_wlast                                 : std_logic;                     -- hps_system:h2f_lw_WLAST -> mm_interconnect_0:hps_system_h2f_lw_axi_master_wlast
	signal hps_system_h2f_lw_axi_master_rresp                                 : std_logic_vector(1 downto 0);  -- mm_interconnect_0:hps_system_h2f_lw_axi_master_rresp -> hps_system:h2f_lw_RRESP
	signal hps_system_h2f_lw_axi_master_awid                                  : std_logic_vector(11 downto 0); -- hps_system:h2f_lw_AWID -> mm_interconnect_0:hps_system_h2f_lw_axi_master_awid
	signal hps_system_h2f_lw_axi_master_bid                                   : std_logic_vector(11 downto 0); -- mm_interconnect_0:hps_system_h2f_lw_axi_master_bid -> hps_system:h2f_lw_BID
	signal hps_system_h2f_lw_axi_master_bvalid                                : std_logic;                     -- mm_interconnect_0:hps_system_h2f_lw_axi_master_bvalid -> hps_system:h2f_lw_BVALID
	signal hps_system_h2f_lw_axi_master_awsize                                : std_logic_vector(2 downto 0);  -- hps_system:h2f_lw_AWSIZE -> mm_interconnect_0:hps_system_h2f_lw_axi_master_awsize
	signal hps_system_h2f_lw_axi_master_awvalid                               : std_logic;                     -- hps_system:h2f_lw_AWVALID -> mm_interconnect_0:hps_system_h2f_lw_axi_master_awvalid
	signal hps_system_h2f_lw_axi_master_rvalid                                : std_logic;                     -- mm_interconnect_0:hps_system_h2f_lw_axi_master_rvalid -> hps_system:h2f_lw_RVALID
	signal master_jtag_master_readdata                                        : std_logic_vector(31 downto 0); -- mm_interconnect_0:master_jtag_master_readdata -> master_jtag:master_readdata
	signal master_jtag_master_waitrequest                                     : std_logic;                     -- mm_interconnect_0:master_jtag_master_waitrequest -> master_jtag:master_waitrequest
	signal master_jtag_master_address                                         : std_logic_vector(31 downto 0); -- master_jtag:master_address -> mm_interconnect_0:master_jtag_master_address
	signal master_jtag_master_read                                            : std_logic;                     -- master_jtag:master_read -> mm_interconnect_0:master_jtag_master_read
	signal master_jtag_master_byteenable                                      : std_logic_vector(3 downto 0);  -- master_jtag:master_byteenable -> mm_interconnect_0:master_jtag_master_byteenable
	signal master_jtag_master_readdatavalid                                   : std_logic;                     -- mm_interconnect_0:master_jtag_master_readdatavalid -> master_jtag:master_readdatavalid
	signal master_jtag_master_write                                           : std_logic;                     -- master_jtag:master_write -> mm_interconnect_0:master_jtag_master_write
	signal master_jtag_master_writedata                                       : std_logic_vector(31 downto 0); -- master_jtag:master_writedata -> mm_interconnect_0:master_jtag_master_writedata
	signal mm_interconnect_0_a_4_quadrant_chopper_0_avalon_slave_0_readdata   : std_logic_vector(15 downto 0); -- a_4_quadrant_chopper_0:avs_readdata -> mm_interconnect_0:a_4_quadrant_chopper_0_avalon_slave_0_readdata
	signal mm_interconnect_0_a_4_quadrant_chopper_0_avalon_slave_0_address    : std_logic_vector(1 downto 0);  -- mm_interconnect_0:a_4_quadrant_chopper_0_avalon_slave_0_address -> a_4_quadrant_chopper_0:avs_address
	signal mm_interconnect_0_a_4_quadrant_chopper_0_avalon_slave_0_read       : std_logic;                     -- mm_interconnect_0:a_4_quadrant_chopper_0_avalon_slave_0_read -> a_4_quadrant_chopper_0:avs_read
	signal mm_interconnect_0_a_4_quadrant_chopper_0_avalon_slave_0_byteenable : std_logic_vector(1 downto 0);  -- mm_interconnect_0:a_4_quadrant_chopper_0_avalon_slave_0_byteenable -> a_4_quadrant_chopper_0:avs_byteenable
	signal mm_interconnect_0_a_4_quadrant_chopper_0_avalon_slave_0_write      : std_logic;                     -- mm_interconnect_0:a_4_quadrant_chopper_0_avalon_slave_0_write -> a_4_quadrant_chopper_0:avs_write
	signal mm_interconnect_0_a_4_quadrant_chopper_0_avalon_slave_0_writedata  : std_logic_vector(15 downto 0); -- mm_interconnect_0:a_4_quadrant_chopper_0_avalon_slave_0_writedata -> a_4_quadrant_chopper_0:avs_writedata
	signal mm_interconnect_0_sysid_control_slave_readdata                     : std_logic_vector(31 downto 0); -- sysid:readdata -> mm_interconnect_0:sysid_control_slave_readdata
	signal mm_interconnect_0_sysid_control_slave_address                      : std_logic_vector(0 downto 0);  -- mm_interconnect_0:sysid_control_slave_address -> sysid:address
	signal a_4_quadrant_chopper_0_interrupt_sender_0_irq                      : std_logic;                     -- a_4_quadrant_chopper_0:ins_end_cycle -> a_4_quadrant_chopper_0_interrupt_sender_0_irq:in
	signal hps_system_f2h_irq0_irq                                            : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> hps_system:f2h_irq_p0
	signal hps_system_f2h_irq1_irq                                            : std_logic_vector(31 downto 0); -- irq_mapper_001:sender_irq -> hps_system:f2h_irq_p1
	signal rst_controller_reset_out_reset                                     : std_logic;                     -- rst_controller:reset_out -> [a_4_quadrant_chopper_0:rsi_reset, mm_interconnect_0:a_4_quadrant_chopper_0_clock_reset_reset_bridge_in_reset_reset, mm_interconnect_0:master_jtag_clk_reset_reset_bridge_in_reset_reset, rst_controller_reset_out_reset:in]
	signal rst_controller_001_reset_out_reset                                 : std_logic;                     -- rst_controller_001:reset_out -> mm_interconnect_0:hps_system_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset
	signal hps_system_h2f_reset_reset                                         : std_logic;                     -- hps_system:h2f_rst_n -> hps_system_h2f_reset_reset:in
	signal reset_reset_n_ports_inv                                            : std_logic;                     -- reset_reset_n:inv -> [master_jtag:clk_reset_reset, rst_controller:reset_in0]
	signal irq_mapper_receiver0_inv                                           : std_logic;                     -- a_4_quadrant_chopper_0_interrupt_sender_0_irq:inv -> irq_mapper:receiver0_irq
	signal rst_controller_reset_out_reset_ports_inv                           : std_logic;                     -- rst_controller_reset_out_reset:inv -> sysid:reset_n
	signal hps_system_h2f_reset_reset_ports_inv                               : std_logic;                     -- hps_system_h2f_reset_reset:inv -> rst_controller_001:reset_in0

begin

	a_4_quadrant_chopper_0 : component hacheur_top
		port map (
			rsi_reset      => rst_controller_reset_out_reset,                                     --        clock_reset.reset
			avs_address    => mm_interconnect_0_a_4_quadrant_chopper_0_avalon_slave_0_address,    --     avalon_slave_0.address
			avs_byteenable => mm_interconnect_0_a_4_quadrant_chopper_0_avalon_slave_0_byteenable, --                   .byteenable
			avs_read       => mm_interconnect_0_a_4_quadrant_chopper_0_avalon_slave_0_read,       --                   .read
			avs_readdata   => mm_interconnect_0_a_4_quadrant_chopper_0_avalon_slave_0_readdata,   --                   .readdata
			avs_write      => mm_interconnect_0_a_4_quadrant_chopper_0_avalon_slave_0_write,      --                   .write
			avs_writedata  => mm_interconnect_0_a_4_quadrant_chopper_0_avalon_slave_0_writedata,  --                   .writedata
			ins_end_cycle  => a_4_quadrant_chopper_0_interrupt_sender_0_irq,                      -- interrupt_sender_0.irq_n
			csi_clock      => clk_clk,                                                            --         clock_sink.clk
			A              => pwm_a_pwm,                                                          --        conduit_end.a_pwm
			B              => pwm_b_pwm,                                                          --                   .b_pwm
			secure         => pwm_secure                                                          --                   .secure
		);

	hps_system : component core_hps_system
		generic map (
			F2S_Width => 2,
			S2F_Width => 2
		)
		port map (
			h2f_mpu_eventi           => open,                                 --    h2f_mpu_events.eventi
			h2f_mpu_evento           => open,                                 --                  .evento
			h2f_mpu_standbywfe       => open,                                 --                  .standbywfe
			h2f_mpu_standbywfi       => open,                                 --                  .standbywfi
			mem_a                    => memory_mem_a,                         --            memory.mem_a
			mem_ba                   => memory_mem_ba,                        --                  .mem_ba
			mem_ck                   => memory_mem_ck,                        --                  .mem_ck
			mem_ck_n                 => memory_mem_ck_n,                      --                  .mem_ck_n
			mem_cke                  => memory_mem_cke,                       --                  .mem_cke
			mem_cs_n                 => memory_mem_cs_n,                      --                  .mem_cs_n
			mem_ras_n                => memory_mem_ras_n,                     --                  .mem_ras_n
			mem_cas_n                => memory_mem_cas_n,                     --                  .mem_cas_n
			mem_we_n                 => memory_mem_we_n,                      --                  .mem_we_n
			mem_reset_n              => memory_mem_reset_n,                   --                  .mem_reset_n
			mem_dq                   => memory_mem_dq,                        --                  .mem_dq
			mem_dqs                  => memory_mem_dqs,                       --                  .mem_dqs
			mem_dqs_n                => memory_mem_dqs_n,                     --                  .mem_dqs_n
			mem_odt                  => memory_mem_odt,                       --                  .mem_odt
			mem_dm                   => memory_mem_dm,                        --                  .mem_dm
			oct_rzqin                => memory_oct_rzqin,                     --                  .oct_rzqin
			hps_io_emac1_inst_TX_CLK => hps_io_hps_io_emac1_inst_TX_CLK,      --            hps_io.hps_io_emac1_inst_TX_CLK
			hps_io_emac1_inst_TXD0   => hps_io_hps_io_emac1_inst_TXD0,        --                  .hps_io_emac1_inst_TXD0
			hps_io_emac1_inst_TXD1   => hps_io_hps_io_emac1_inst_TXD1,        --                  .hps_io_emac1_inst_TXD1
			hps_io_emac1_inst_TXD2   => hps_io_hps_io_emac1_inst_TXD2,        --                  .hps_io_emac1_inst_TXD2
			hps_io_emac1_inst_TXD3   => hps_io_hps_io_emac1_inst_TXD3,        --                  .hps_io_emac1_inst_TXD3
			hps_io_emac1_inst_RXD0   => hps_io_hps_io_emac1_inst_RXD0,        --                  .hps_io_emac1_inst_RXD0
			hps_io_emac1_inst_MDIO   => hps_io_hps_io_emac1_inst_MDIO,        --                  .hps_io_emac1_inst_MDIO
			hps_io_emac1_inst_MDC    => hps_io_hps_io_emac1_inst_MDC,         --                  .hps_io_emac1_inst_MDC
			hps_io_emac1_inst_RX_CTL => hps_io_hps_io_emac1_inst_RX_CTL,      --                  .hps_io_emac1_inst_RX_CTL
			hps_io_emac1_inst_TX_CTL => hps_io_hps_io_emac1_inst_TX_CTL,      --                  .hps_io_emac1_inst_TX_CTL
			hps_io_emac1_inst_RX_CLK => hps_io_hps_io_emac1_inst_RX_CLK,      --                  .hps_io_emac1_inst_RX_CLK
			hps_io_emac1_inst_RXD1   => hps_io_hps_io_emac1_inst_RXD1,        --                  .hps_io_emac1_inst_RXD1
			hps_io_emac1_inst_RXD2   => hps_io_hps_io_emac1_inst_RXD2,        --                  .hps_io_emac1_inst_RXD2
			hps_io_emac1_inst_RXD3   => hps_io_hps_io_emac1_inst_RXD3,        --                  .hps_io_emac1_inst_RXD3
			hps_io_sdio_inst_CMD     => hps_io_hps_io_sdio_inst_CMD,          --                  .hps_io_sdio_inst_CMD
			hps_io_sdio_inst_D0      => hps_io_hps_io_sdio_inst_D0,           --                  .hps_io_sdio_inst_D0
			hps_io_sdio_inst_D1      => hps_io_hps_io_sdio_inst_D1,           --                  .hps_io_sdio_inst_D1
			hps_io_sdio_inst_CLK     => hps_io_hps_io_sdio_inst_CLK,          --                  .hps_io_sdio_inst_CLK
			hps_io_sdio_inst_D2      => hps_io_hps_io_sdio_inst_D2,           --                  .hps_io_sdio_inst_D2
			hps_io_sdio_inst_D3      => hps_io_hps_io_sdio_inst_D3,           --                  .hps_io_sdio_inst_D3
			hps_io_uart0_inst_RX     => hps_io_hps_io_uart0_inst_RX,          --                  .hps_io_uart0_inst_RX
			hps_io_uart0_inst_TX     => hps_io_hps_io_uart0_inst_TX,          --                  .hps_io_uart0_inst_TX
			hps_io_i2c0_inst_SDA     => hps_io_hps_io_i2c0_inst_SDA,          --                  .hps_io_i2c0_inst_SDA
			hps_io_i2c0_inst_SCL     => hps_io_hps_io_i2c0_inst_SCL,          --                  .hps_io_i2c0_inst_SCL
			hps_io_i2c1_inst_SDA     => hps_io_hps_io_i2c1_inst_SDA,          --                  .hps_io_i2c1_inst_SDA
			hps_io_i2c1_inst_SCL     => hps_io_hps_io_i2c1_inst_SCL,          --                  .hps_io_i2c1_inst_SCL
			h2f_rst_n                => hps_system_h2f_reset_reset,           --         h2f_reset.reset_n
			f2h_sdram0_clk           => clk_clk,                              --  f2h_sdram0_clock.clk
			f2h_sdram0_ARADDR        => open,                                 --   f2h_sdram0_data.araddr
			f2h_sdram0_ARLEN         => open,                                 --                  .arlen
			f2h_sdram0_ARID          => open,                                 --                  .arid
			f2h_sdram0_ARSIZE        => open,                                 --                  .arsize
			f2h_sdram0_ARBURST       => open,                                 --                  .arburst
			f2h_sdram0_ARLOCK        => open,                                 --                  .arlock
			f2h_sdram0_ARPROT        => open,                                 --                  .arprot
			f2h_sdram0_ARVALID       => open,                                 --                  .arvalid
			f2h_sdram0_ARCACHE       => open,                                 --                  .arcache
			f2h_sdram0_AWADDR        => open,                                 --                  .awaddr
			f2h_sdram0_AWLEN         => open,                                 --                  .awlen
			f2h_sdram0_AWID          => open,                                 --                  .awid
			f2h_sdram0_AWSIZE        => open,                                 --                  .awsize
			f2h_sdram0_AWBURST       => open,                                 --                  .awburst
			f2h_sdram0_AWLOCK        => open,                                 --                  .awlock
			f2h_sdram0_AWPROT        => open,                                 --                  .awprot
			f2h_sdram0_AWVALID       => open,                                 --                  .awvalid
			f2h_sdram0_AWCACHE       => open,                                 --                  .awcache
			f2h_sdram0_BRESP         => open,                                 --                  .bresp
			f2h_sdram0_BID           => open,                                 --                  .bid
			f2h_sdram0_BVALID        => open,                                 --                  .bvalid
			f2h_sdram0_BREADY        => open,                                 --                  .bready
			f2h_sdram0_ARREADY       => open,                                 --                  .arready
			f2h_sdram0_AWREADY       => open,                                 --                  .awready
			f2h_sdram0_RREADY        => open,                                 --                  .rready
			f2h_sdram0_RDATA         => open,                                 --                  .rdata
			f2h_sdram0_RRESP         => open,                                 --                  .rresp
			f2h_sdram0_RLAST         => open,                                 --                  .rlast
			f2h_sdram0_RID           => open,                                 --                  .rid
			f2h_sdram0_RVALID        => open,                                 --                  .rvalid
			f2h_sdram0_WLAST         => open,                                 --                  .wlast
			f2h_sdram0_WVALID        => open,                                 --                  .wvalid
			f2h_sdram0_WDATA         => open,                                 --                  .wdata
			f2h_sdram0_WSTRB         => open,                                 --                  .wstrb
			f2h_sdram0_WREADY        => open,                                 --                  .wready
			f2h_sdram0_WID           => open,                                 --                  .wid
			h2f_axi_clk              => clk_clk,                              --     h2f_axi_clock.clk
			h2f_AWID                 => open,                                 --    h2f_axi_master.awid
			h2f_AWADDR               => open,                                 --                  .awaddr
			h2f_AWLEN                => open,                                 --                  .awlen
			h2f_AWSIZE               => open,                                 --                  .awsize
			h2f_AWBURST              => open,                                 --                  .awburst
			h2f_AWLOCK               => open,                                 --                  .awlock
			h2f_AWCACHE              => open,                                 --                  .awcache
			h2f_AWPROT               => open,                                 --                  .awprot
			h2f_AWVALID              => open,                                 --                  .awvalid
			h2f_AWREADY              => open,                                 --                  .awready
			h2f_WID                  => open,                                 --                  .wid
			h2f_WDATA                => open,                                 --                  .wdata
			h2f_WSTRB                => open,                                 --                  .wstrb
			h2f_WLAST                => open,                                 --                  .wlast
			h2f_WVALID               => open,                                 --                  .wvalid
			h2f_WREADY               => open,                                 --                  .wready
			h2f_BID                  => open,                                 --                  .bid
			h2f_BRESP                => open,                                 --                  .bresp
			h2f_BVALID               => open,                                 --                  .bvalid
			h2f_BREADY               => open,                                 --                  .bready
			h2f_ARID                 => open,                                 --                  .arid
			h2f_ARADDR               => open,                                 --                  .araddr
			h2f_ARLEN                => open,                                 --                  .arlen
			h2f_ARSIZE               => open,                                 --                  .arsize
			h2f_ARBURST              => open,                                 --                  .arburst
			h2f_ARLOCK               => open,                                 --                  .arlock
			h2f_ARCACHE              => open,                                 --                  .arcache
			h2f_ARPROT               => open,                                 --                  .arprot
			h2f_ARVALID              => open,                                 --                  .arvalid
			h2f_ARREADY              => open,                                 --                  .arready
			h2f_RID                  => open,                                 --                  .rid
			h2f_RDATA                => open,                                 --                  .rdata
			h2f_RRESP                => open,                                 --                  .rresp
			h2f_RLAST                => open,                                 --                  .rlast
			h2f_RVALID               => open,                                 --                  .rvalid
			h2f_RREADY               => open,                                 --                  .rready
			f2h_axi_clk              => clk_clk,                              --     f2h_axi_clock.clk
			f2h_AWID                 => open,                                 --     f2h_axi_slave.awid
			f2h_AWADDR               => open,                                 --                  .awaddr
			f2h_AWLEN                => open,                                 --                  .awlen
			f2h_AWSIZE               => open,                                 --                  .awsize
			f2h_AWBURST              => open,                                 --                  .awburst
			f2h_AWLOCK               => open,                                 --                  .awlock
			f2h_AWCACHE              => open,                                 --                  .awcache
			f2h_AWPROT               => open,                                 --                  .awprot
			f2h_AWVALID              => open,                                 --                  .awvalid
			f2h_AWREADY              => open,                                 --                  .awready
			f2h_AWUSER               => open,                                 --                  .awuser
			f2h_WID                  => open,                                 --                  .wid
			f2h_WDATA                => open,                                 --                  .wdata
			f2h_WSTRB                => open,                                 --                  .wstrb
			f2h_WLAST                => open,                                 --                  .wlast
			f2h_WVALID               => open,                                 --                  .wvalid
			f2h_WREADY               => open,                                 --                  .wready
			f2h_BID                  => open,                                 --                  .bid
			f2h_BRESP                => open,                                 --                  .bresp
			f2h_BVALID               => open,                                 --                  .bvalid
			f2h_BREADY               => open,                                 --                  .bready
			f2h_ARID                 => open,                                 --                  .arid
			f2h_ARADDR               => open,                                 --                  .araddr
			f2h_ARLEN                => open,                                 --                  .arlen
			f2h_ARSIZE               => open,                                 --                  .arsize
			f2h_ARBURST              => open,                                 --                  .arburst
			f2h_ARLOCK               => open,                                 --                  .arlock
			f2h_ARCACHE              => open,                                 --                  .arcache
			f2h_ARPROT               => open,                                 --                  .arprot
			f2h_ARVALID              => open,                                 --                  .arvalid
			f2h_ARREADY              => open,                                 --                  .arready
			f2h_ARUSER               => open,                                 --                  .aruser
			f2h_RID                  => open,                                 --                  .rid
			f2h_RDATA                => open,                                 --                  .rdata
			f2h_RRESP                => open,                                 --                  .rresp
			f2h_RLAST                => open,                                 --                  .rlast
			f2h_RVALID               => open,                                 --                  .rvalid
			f2h_RREADY               => open,                                 --                  .rready
			h2f_lw_axi_clk           => clk_clk,                              --  h2f_lw_axi_clock.clk
			h2f_lw_AWID              => hps_system_h2f_lw_axi_master_awid,    -- h2f_lw_axi_master.awid
			h2f_lw_AWADDR            => hps_system_h2f_lw_axi_master_awaddr,  --                  .awaddr
			h2f_lw_AWLEN             => hps_system_h2f_lw_axi_master_awlen,   --                  .awlen
			h2f_lw_AWSIZE            => hps_system_h2f_lw_axi_master_awsize,  --                  .awsize
			h2f_lw_AWBURST           => hps_system_h2f_lw_axi_master_awburst, --                  .awburst
			h2f_lw_AWLOCK            => hps_system_h2f_lw_axi_master_awlock,  --                  .awlock
			h2f_lw_AWCACHE           => hps_system_h2f_lw_axi_master_awcache, --                  .awcache
			h2f_lw_AWPROT            => hps_system_h2f_lw_axi_master_awprot,  --                  .awprot
			h2f_lw_AWVALID           => hps_system_h2f_lw_axi_master_awvalid, --                  .awvalid
			h2f_lw_AWREADY           => hps_system_h2f_lw_axi_master_awready, --                  .awready
			h2f_lw_WID               => hps_system_h2f_lw_axi_master_wid,     --                  .wid
			h2f_lw_WDATA             => hps_system_h2f_lw_axi_master_wdata,   --                  .wdata
			h2f_lw_WSTRB             => hps_system_h2f_lw_axi_master_wstrb,   --                  .wstrb
			h2f_lw_WLAST             => hps_system_h2f_lw_axi_master_wlast,   --                  .wlast
			h2f_lw_WVALID            => hps_system_h2f_lw_axi_master_wvalid,  --                  .wvalid
			h2f_lw_WREADY            => hps_system_h2f_lw_axi_master_wready,  --                  .wready
			h2f_lw_BID               => hps_system_h2f_lw_axi_master_bid,     --                  .bid
			h2f_lw_BRESP             => hps_system_h2f_lw_axi_master_bresp,   --                  .bresp
			h2f_lw_BVALID            => hps_system_h2f_lw_axi_master_bvalid,  --                  .bvalid
			h2f_lw_BREADY            => hps_system_h2f_lw_axi_master_bready,  --                  .bready
			h2f_lw_ARID              => hps_system_h2f_lw_axi_master_arid,    --                  .arid
			h2f_lw_ARADDR            => hps_system_h2f_lw_axi_master_araddr,  --                  .araddr
			h2f_lw_ARLEN             => hps_system_h2f_lw_axi_master_arlen,   --                  .arlen
			h2f_lw_ARSIZE            => hps_system_h2f_lw_axi_master_arsize,  --                  .arsize
			h2f_lw_ARBURST           => hps_system_h2f_lw_axi_master_arburst, --                  .arburst
			h2f_lw_ARLOCK            => hps_system_h2f_lw_axi_master_arlock,  --                  .arlock
			h2f_lw_ARCACHE           => hps_system_h2f_lw_axi_master_arcache, --                  .arcache
			h2f_lw_ARPROT            => hps_system_h2f_lw_axi_master_arprot,  --                  .arprot
			h2f_lw_ARVALID           => hps_system_h2f_lw_axi_master_arvalid, --                  .arvalid
			h2f_lw_ARREADY           => hps_system_h2f_lw_axi_master_arready, --                  .arready
			h2f_lw_RID               => hps_system_h2f_lw_axi_master_rid,     --                  .rid
			h2f_lw_RDATA             => hps_system_h2f_lw_axi_master_rdata,   --                  .rdata
			h2f_lw_RRESP             => hps_system_h2f_lw_axi_master_rresp,   --                  .rresp
			h2f_lw_RLAST             => hps_system_h2f_lw_axi_master_rlast,   --                  .rlast
			h2f_lw_RVALID            => hps_system_h2f_lw_axi_master_rvalid,  --                  .rvalid
			h2f_lw_RREADY            => hps_system_h2f_lw_axi_master_rready,  --                  .rready
			f2h_irq_p0               => hps_system_f2h_irq0_irq,              --          f2h_irq0.irq
			f2h_irq_p1               => hps_system_f2h_irq1_irq               --          f2h_irq1.irq
		);

	master_jtag : component core_master_jtag
		generic map (
			USE_PLI     => 0,
			PLI_PORT    => 50000,
			FIFO_DEPTHS => 2
		)
		port map (
			clk_clk              => clk_clk,                          --          clk.clk
			clk_reset_reset      => reset_reset_n_ports_inv,          --    clk_reset.reset
			master_address       => master_jtag_master_address,       --       master.address
			master_readdata      => master_jtag_master_readdata,      --             .readdata
			master_read          => master_jtag_master_read,          --             .read
			master_write         => master_jtag_master_write,         --             .write
			master_writedata     => master_jtag_master_writedata,     --             .writedata
			master_waitrequest   => master_jtag_master_waitrequest,   --             .waitrequest
			master_readdatavalid => master_jtag_master_readdatavalid, --             .readdatavalid
			master_byteenable    => master_jtag_master_byteenable,    --             .byteenable
			master_reset_reset   => open                              -- master_reset.reset
		);

	sysid : component core_sysid
		port map (
			clock    => clk_clk,                                          --           clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,         --         reset.reset_n
			readdata => mm_interconnect_0_sysid_control_slave_readdata,   -- control_slave.readdata
			address  => mm_interconnect_0_sysid_control_slave_address(0)  --              .address
		);

	mm_interconnect_0 : component core_mm_interconnect_0
		port map (
			hps_system_h2f_lw_axi_master_awid                                        => hps_system_h2f_lw_axi_master_awid,                                  --                                       hps_system_h2f_lw_axi_master.awid
			hps_system_h2f_lw_axi_master_awaddr                                      => hps_system_h2f_lw_axi_master_awaddr,                                --                                                                   .awaddr
			hps_system_h2f_lw_axi_master_awlen                                       => hps_system_h2f_lw_axi_master_awlen,                                 --                                                                   .awlen
			hps_system_h2f_lw_axi_master_awsize                                      => hps_system_h2f_lw_axi_master_awsize,                                --                                                                   .awsize
			hps_system_h2f_lw_axi_master_awburst                                     => hps_system_h2f_lw_axi_master_awburst,                               --                                                                   .awburst
			hps_system_h2f_lw_axi_master_awlock                                      => hps_system_h2f_lw_axi_master_awlock,                                --                                                                   .awlock
			hps_system_h2f_lw_axi_master_awcache                                     => hps_system_h2f_lw_axi_master_awcache,                               --                                                                   .awcache
			hps_system_h2f_lw_axi_master_awprot                                      => hps_system_h2f_lw_axi_master_awprot,                                --                                                                   .awprot
			hps_system_h2f_lw_axi_master_awvalid                                     => hps_system_h2f_lw_axi_master_awvalid,                               --                                                                   .awvalid
			hps_system_h2f_lw_axi_master_awready                                     => hps_system_h2f_lw_axi_master_awready,                               --                                                                   .awready
			hps_system_h2f_lw_axi_master_wid                                         => hps_system_h2f_lw_axi_master_wid,                                   --                                                                   .wid
			hps_system_h2f_lw_axi_master_wdata                                       => hps_system_h2f_lw_axi_master_wdata,                                 --                                                                   .wdata
			hps_system_h2f_lw_axi_master_wstrb                                       => hps_system_h2f_lw_axi_master_wstrb,                                 --                                                                   .wstrb
			hps_system_h2f_lw_axi_master_wlast                                       => hps_system_h2f_lw_axi_master_wlast,                                 --                                                                   .wlast
			hps_system_h2f_lw_axi_master_wvalid                                      => hps_system_h2f_lw_axi_master_wvalid,                                --                                                                   .wvalid
			hps_system_h2f_lw_axi_master_wready                                      => hps_system_h2f_lw_axi_master_wready,                                --                                                                   .wready
			hps_system_h2f_lw_axi_master_bid                                         => hps_system_h2f_lw_axi_master_bid,                                   --                                                                   .bid
			hps_system_h2f_lw_axi_master_bresp                                       => hps_system_h2f_lw_axi_master_bresp,                                 --                                                                   .bresp
			hps_system_h2f_lw_axi_master_bvalid                                      => hps_system_h2f_lw_axi_master_bvalid,                                --                                                                   .bvalid
			hps_system_h2f_lw_axi_master_bready                                      => hps_system_h2f_lw_axi_master_bready,                                --                                                                   .bready
			hps_system_h2f_lw_axi_master_arid                                        => hps_system_h2f_lw_axi_master_arid,                                  --                                                                   .arid
			hps_system_h2f_lw_axi_master_araddr                                      => hps_system_h2f_lw_axi_master_araddr,                                --                                                                   .araddr
			hps_system_h2f_lw_axi_master_arlen                                       => hps_system_h2f_lw_axi_master_arlen,                                 --                                                                   .arlen
			hps_system_h2f_lw_axi_master_arsize                                      => hps_system_h2f_lw_axi_master_arsize,                                --                                                                   .arsize
			hps_system_h2f_lw_axi_master_arburst                                     => hps_system_h2f_lw_axi_master_arburst,                               --                                                                   .arburst
			hps_system_h2f_lw_axi_master_arlock                                      => hps_system_h2f_lw_axi_master_arlock,                                --                                                                   .arlock
			hps_system_h2f_lw_axi_master_arcache                                     => hps_system_h2f_lw_axi_master_arcache,                               --                                                                   .arcache
			hps_system_h2f_lw_axi_master_arprot                                      => hps_system_h2f_lw_axi_master_arprot,                                --                                                                   .arprot
			hps_system_h2f_lw_axi_master_arvalid                                     => hps_system_h2f_lw_axi_master_arvalid,                               --                                                                   .arvalid
			hps_system_h2f_lw_axi_master_arready                                     => hps_system_h2f_lw_axi_master_arready,                               --                                                                   .arready
			hps_system_h2f_lw_axi_master_rid                                         => hps_system_h2f_lw_axi_master_rid,                                   --                                                                   .rid
			hps_system_h2f_lw_axi_master_rdata                                       => hps_system_h2f_lw_axi_master_rdata,                                 --                                                                   .rdata
			hps_system_h2f_lw_axi_master_rresp                                       => hps_system_h2f_lw_axi_master_rresp,                                 --                                                                   .rresp
			hps_system_h2f_lw_axi_master_rlast                                       => hps_system_h2f_lw_axi_master_rlast,                                 --                                                                   .rlast
			hps_system_h2f_lw_axi_master_rvalid                                      => hps_system_h2f_lw_axi_master_rvalid,                                --                                                                   .rvalid
			hps_system_h2f_lw_axi_master_rready                                      => hps_system_h2f_lw_axi_master_rready,                                --                                                                   .rready
			clk_0_clk_clk                                                            => clk_clk,                                                            --                                                          clk_0_clk.clk
			a_4_quadrant_chopper_0_clock_reset_reset_bridge_in_reset_reset           => rst_controller_reset_out_reset,                                     --           a_4_quadrant_chopper_0_clock_reset_reset_bridge_in_reset.reset
			hps_system_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset => rst_controller_001_reset_out_reset,                                 -- hps_system_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
			master_jtag_clk_reset_reset_bridge_in_reset_reset                        => rst_controller_reset_out_reset,                                     --                        master_jtag_clk_reset_reset_bridge_in_reset.reset
			master_jtag_master_address                                               => master_jtag_master_address,                                         --                                                 master_jtag_master.address
			master_jtag_master_waitrequest                                           => master_jtag_master_waitrequest,                                     --                                                                   .waitrequest
			master_jtag_master_byteenable                                            => master_jtag_master_byteenable,                                      --                                                                   .byteenable
			master_jtag_master_read                                                  => master_jtag_master_read,                                            --                                                                   .read
			master_jtag_master_readdata                                              => master_jtag_master_readdata,                                        --                                                                   .readdata
			master_jtag_master_readdatavalid                                         => master_jtag_master_readdatavalid,                                   --                                                                   .readdatavalid
			master_jtag_master_write                                                 => master_jtag_master_write,                                           --                                                                   .write
			master_jtag_master_writedata                                             => master_jtag_master_writedata,                                       --                                                                   .writedata
			a_4_quadrant_chopper_0_avalon_slave_0_address                            => mm_interconnect_0_a_4_quadrant_chopper_0_avalon_slave_0_address,    --                              a_4_quadrant_chopper_0_avalon_slave_0.address
			a_4_quadrant_chopper_0_avalon_slave_0_write                              => mm_interconnect_0_a_4_quadrant_chopper_0_avalon_slave_0_write,      --                                                                   .write
			a_4_quadrant_chopper_0_avalon_slave_0_read                               => mm_interconnect_0_a_4_quadrant_chopper_0_avalon_slave_0_read,       --                                                                   .read
			a_4_quadrant_chopper_0_avalon_slave_0_readdata                           => mm_interconnect_0_a_4_quadrant_chopper_0_avalon_slave_0_readdata,   --                                                                   .readdata
			a_4_quadrant_chopper_0_avalon_slave_0_writedata                          => mm_interconnect_0_a_4_quadrant_chopper_0_avalon_slave_0_writedata,  --                                                                   .writedata
			a_4_quadrant_chopper_0_avalon_slave_0_byteenable                         => mm_interconnect_0_a_4_quadrant_chopper_0_avalon_slave_0_byteenable, --                                                                   .byteenable
			sysid_control_slave_address                                              => mm_interconnect_0_sysid_control_slave_address,                      --                                                sysid_control_slave.address
			sysid_control_slave_readdata                                             => mm_interconnect_0_sysid_control_slave_readdata                      --                                                                   .readdata
		);

	irq_mapper : component core_irq_mapper
		port map (
			clk           => open,                     --       clk.clk
			reset         => open,                     -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_inv, -- receiver0.irq
			sender_irq    => hps_system_f2h_irq0_irq   --    sender.irq
		);

	irq_mapper_001 : component core_irq_mapper_001
		port map (
			clk        => open,                    --       clk.clk
			reset      => open,                    -- clk_reset.reset
			sender_irq => hps_system_f2h_irq1_irq  --    sender.irq
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,        -- reset_in0.reset
			clk            => clk_clk,                        --       clk.clk
			reset_out      => rst_controller_reset_out_reset, -- reset_out.reset
			reset_req      => open,                           -- (terminated)
			reset_req_in0  => '0',                            -- (terminated)
			reset_in1      => '0',                            -- (terminated)
			reset_req_in1  => '0',                            -- (terminated)
			reset_in2      => '0',                            -- (terminated)
			reset_req_in2  => '0',                            -- (terminated)
			reset_in3      => '0',                            -- (terminated)
			reset_req_in3  => '0',                            -- (terminated)
			reset_in4      => '0',                            -- (terminated)
			reset_req_in4  => '0',                            -- (terminated)
			reset_in5      => '0',                            -- (terminated)
			reset_req_in5  => '0',                            -- (terminated)
			reset_in6      => '0',                            -- (terminated)
			reset_req_in6  => '0',                            -- (terminated)
			reset_in7      => '0',                            -- (terminated)
			reset_req_in7  => '0',                            -- (terminated)
			reset_in8      => '0',                            -- (terminated)
			reset_req_in8  => '0',                            -- (terminated)
			reset_in9      => '0',                            -- (terminated)
			reset_req_in9  => '0',                            -- (terminated)
			reset_in10     => '0',                            -- (terminated)
			reset_req_in10 => '0',                            -- (terminated)
			reset_in11     => '0',                            -- (terminated)
			reset_req_in11 => '0',                            -- (terminated)
			reset_in12     => '0',                            -- (terminated)
			reset_req_in12 => '0',                            -- (terminated)
			reset_in13     => '0',                            -- (terminated)
			reset_req_in13 => '0',                            -- (terminated)
			reset_in14     => '0',                            -- (terminated)
			reset_req_in14 => '0',                            -- (terminated)
			reset_in15     => '0',                            -- (terminated)
			reset_req_in15 => '0'                             -- (terminated)
		);

	rst_controller_001 : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => hps_system_h2f_reset_reset_ports_inv, -- reset_in0.reset
			clk            => clk_clk,                              --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset,   -- reset_out.reset
			reset_req      => open,                                 -- (terminated)
			reset_req_in0  => '0',                                  -- (terminated)
			reset_in1      => '0',                                  -- (terminated)
			reset_req_in1  => '0',                                  -- (terminated)
			reset_in2      => '0',                                  -- (terminated)
			reset_req_in2  => '0',                                  -- (terminated)
			reset_in3      => '0',                                  -- (terminated)
			reset_req_in3  => '0',                                  -- (terminated)
			reset_in4      => '0',                                  -- (terminated)
			reset_req_in4  => '0',                                  -- (terminated)
			reset_in5      => '0',                                  -- (terminated)
			reset_req_in5  => '0',                                  -- (terminated)
			reset_in6      => '0',                                  -- (terminated)
			reset_req_in6  => '0',                                  -- (terminated)
			reset_in7      => '0',                                  -- (terminated)
			reset_req_in7  => '0',                                  -- (terminated)
			reset_in8      => '0',                                  -- (terminated)
			reset_req_in8  => '0',                                  -- (terminated)
			reset_in9      => '0',                                  -- (terminated)
			reset_req_in9  => '0',                                  -- (terminated)
			reset_in10     => '0',                                  -- (terminated)
			reset_req_in10 => '0',                                  -- (terminated)
			reset_in11     => '0',                                  -- (terminated)
			reset_req_in11 => '0',                                  -- (terminated)
			reset_in12     => '0',                                  -- (terminated)
			reset_req_in12 => '0',                                  -- (terminated)
			reset_in13     => '0',                                  -- (terminated)
			reset_req_in13 => '0',                                  -- (terminated)
			reset_in14     => '0',                                  -- (terminated)
			reset_req_in14 => '0',                                  -- (terminated)
			reset_in15     => '0',                                  -- (terminated)
			reset_req_in15 => '0'                                   -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	irq_mapper_receiver0_inv <= not a_4_quadrant_chopper_0_interrupt_sender_0_irq;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

	hps_system_h2f_reset_reset_ports_inv <= not hps_system_h2f_reset_reset;

end architecture rtl; -- of core
